VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pwm_top
  CLASS BLOCK ;
  FOREIGN pwm_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2300.000 BY 1000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 10.920 2300.000 11.520 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 677.320 2300.000 677.920 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 743.960 2300.000 744.560 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 810.600 2300.000 811.200 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 877.240 2300.000 877.840 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 943.880 2300.000 944.480 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2256.850 996.000 2257.130 1000.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2001.550 996.000 2001.830 1000.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.790 996.000 1746.070 1000.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.490 996.000 1490.770 1000.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1234.730 996.000 1235.010 1000.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 77.560 2300.000 78.160 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.430 996.000 979.710 1000.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.670 996.000 723.950 1000.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 996.000 468.190 1000.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 996.000 212.890 1000.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 987.400 4.000 988.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 916.000 4.000 916.600 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 844.600 4.000 845.200 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.200 4.000 773.800 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.800 4.000 702.400 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 630.400 4.000 631.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 144.200 2300.000 144.800 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 487.600 4.000 488.200 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.800 4.000 345.400 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 210.840 2300.000 211.440 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 277.480 2300.000 278.080 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 344.120 2300.000 344.720 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 410.760 2300.000 411.360 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 477.400 2300.000 478.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 544.040 2300.000 544.640 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 610.680 2300.000 611.280 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 55.120 2300.000 55.720 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 722.200 2300.000 722.800 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 788.840 2300.000 789.440 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 855.480 2300.000 856.080 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 922.120 2300.000 922.720 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 988.760 2300.000 989.360 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2086.650 996.000 2086.930 1000.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1830.890 996.000 1831.170 1000.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.590 996.000 1575.870 1000.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.830 996.000 1320.110 1000.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.530 996.000 1064.810 1000.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 121.760 2300.000 122.360 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.770 996.000 809.050 1000.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 996.000 553.750 1000.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 996.000 297.990 1000.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 996.000 42.690 1000.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.800 4.000 940.400 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 868.400 4.000 869.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 725.600 4.000 726.200 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.800 4.000 583.400 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 188.400 2300.000 189.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.000 4.000 440.600 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 255.040 2300.000 255.640 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 321.680 2300.000 322.280 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 388.320 2300.000 388.920 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 454.960 2300.000 455.560 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 521.600 2300.000 522.200 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 588.240 2300.000 588.840 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 654.880 2300.000 655.480 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 32.680 2300.000 33.280 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 699.760 2300.000 700.360 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 766.400 2300.000 767.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 833.040 2300.000 833.640 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 899.680 2300.000 900.280 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 966.320 2300.000 966.920 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2171.750 996.000 2172.030 1000.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1916.450 996.000 1916.730 1000.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1660.690 996.000 1660.970 1000.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.930 996.000 1405.210 1000.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 996.000 1149.910 1000.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 99.320 2300.000 99.920 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.870 996.000 894.150 1000.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 996.000 638.850 1000.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 996.000 383.090 1000.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 996.000 127.790 1000.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 963.600 4.000 964.200 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.200 4.000 892.800 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.800 4.000 821.400 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 165.960 2300.000 166.560 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.200 4.000 535.800 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 4.000 393.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 232.600 2300.000 233.200 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 299.240 2300.000 299.840 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 366.560 2300.000 367.160 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 433.200 2300.000 433.800 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 499.840 2300.000 500.440 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 566.480 2300.000 567.080 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2296.000 633.120 2300.000 633.720 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2288.130 0.000 2288.410 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2292.730 0.000 2293.010 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2297.330 0.000 2297.610 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1896.210 0.000 1896.490 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1910.470 0.000 1910.750 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1924.270 0.000 1924.550 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.070 0.000 1938.350 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1952.330 0.000 1952.610 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1966.130 0.000 1966.410 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.390 0.000 1980.670 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.190 0.000 1994.470 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2008.450 0.000 2008.730 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2022.250 0.000 2022.530 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.730 0.000 637.010 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2036.050 0.000 2036.330 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2050.310 0.000 2050.590 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2064.110 0.000 2064.390 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2078.370 0.000 2078.650 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2092.170 0.000 2092.450 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.430 0.000 2106.710 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2120.230 0.000 2120.510 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2134.030 0.000 2134.310 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.290 0.000 2148.570 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2162.090 0.000 2162.370 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2176.350 0.000 2176.630 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2190.150 0.000 2190.430 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2204.410 0.000 2204.690 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.210 0.000 2218.490 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2232.010 0.000 2232.290 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2246.270 0.000 2246.550 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.070 0.000 2260.350 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2274.330 0.000 2274.610 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 0.000 665.070 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 0.000 678.870 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 0.000 693.130 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 0.000 706.930 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 0.000 720.730 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.710 0.000 734.990 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.510 0.000 748.790 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.770 0.000 763.050 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 0.000 776.850 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.370 0.000 790.650 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 0.000 804.910 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 0.000 818.710 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.690 0.000 832.970 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 0.000 846.770 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.750 0.000 861.030 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.550 0.000 874.830 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.350 0.000 888.630 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 0.000 902.890 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.410 0.000 916.690 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.670 0.000 930.950 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.470 0.000 944.750 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.730 0.000 959.010 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 0.000 972.810 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.330 0.000 986.610 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.590 0.000 1000.870 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 0.000 1014.670 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.650 0.000 1028.930 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.450 0.000 1042.730 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 0.000 539.030 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.710 0.000 1056.990 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.510 0.000 1070.790 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.310 0.000 1084.590 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.570 0.000 1098.850 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.370 0.000 1112.650 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.630 0.000 1126.910 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.430 0.000 1140.710 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.690 0.000 1154.970 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.490 0.000 1168.770 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.290 0.000 1182.570 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 0.000 552.830 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.550 0.000 1196.830 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.350 0.000 1210.630 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.610 0.000 1224.890 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.410 0.000 1238.690 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 0.000 1252.950 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.470 0.000 1266.750 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.270 0.000 1280.550 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.530 0.000 1294.810 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.330 0.000 1308.610 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.590 0.000 1322.870 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.390 0.000 1336.670 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.650 0.000 1350.930 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.450 0.000 1364.730 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.250 0.000 1378.530 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.510 0.000 1392.790 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.310 0.000 1406.590 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.570 0.000 1420.850 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1434.370 0.000 1434.650 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1448.630 0.000 1448.910 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.430 0.000 1462.710 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1476.230 0.000 1476.510 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.490 0.000 1490.770 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1504.290 0.000 1504.570 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.550 0.000 1518.830 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.350 0.000 1532.630 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1546.150 0.000 1546.430 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1560.410 0.000 1560.690 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.210 0.000 1574.490 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.470 0.000 1588.750 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1602.270 0.000 1602.550 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 0.000 595.150 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.530 0.000 1616.810 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1630.330 0.000 1630.610 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1644.130 0.000 1644.410 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.390 0.000 1658.670 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.190 0.000 1672.470 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1686.450 0.000 1686.730 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.250 0.000 1700.530 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1714.510 0.000 1714.790 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.310 0.000 1728.590 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.110 0.000 1742.390 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.370 0.000 1756.650 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.170 0.000 1770.450 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1784.430 0.000 1784.710 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1798.230 0.000 1798.510 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.490 0.000 1812.770 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1826.290 0.000 1826.570 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.090 0.000 1840.370 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.350 0.000 1854.630 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.150 0.000 1868.430 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.410 0.000 1882.690 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 0.000 622.750 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 0.000 501.770 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1900.810 0.000 1901.090 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.070 0.000 1915.350 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1928.870 0.000 1929.150 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1943.130 0.000 1943.410 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1956.930 0.000 1957.210 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1970.730 0.000 1971.010 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1984.990 0.000 1985.270 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1998.790 0.000 1999.070 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2013.050 0.000 2013.330 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2026.850 0.000 2027.130 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 0.000 641.610 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.110 0.000 2041.390 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2054.910 0.000 2055.190 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.710 0.000 2068.990 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2082.970 0.000 2083.250 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2096.770 0.000 2097.050 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2111.030 0.000 2111.310 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.830 0.000 2125.110 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2139.090 0.000 2139.370 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2152.890 0.000 2153.170 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.690 0.000 2166.970 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 0.000 655.410 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.950 0.000 2181.230 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2194.750 0.000 2195.030 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2209.010 0.000 2209.290 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2222.810 0.000 2223.090 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2237.070 0.000 2237.350 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2250.870 0.000 2251.150 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2264.670 0.000 2264.950 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.930 0.000 2279.210 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.390 0.000 669.670 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 0.000 683.470 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 0.000 711.530 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.510 0.000 725.790 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 0.000 739.590 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.110 0.000 753.390 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 0.000 781.450 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 0.000 795.710 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.230 0.000 809.510 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.030 0.000 823.310 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 0.000 851.370 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.350 0.000 865.630 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.410 0.000 893.690 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.210 0.000 907.490 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.010 0.000 921.290 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.270 0.000 935.550 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.070 0.000 949.350 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.330 0.000 963.610 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.130 0.000 977.410 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.390 0.000 991.670 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.190 0.000 1005.470 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.990 0.000 1019.270 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.250 0.000 1033.530 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.050 0.000 1047.330 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 0.000 543.630 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.310 0.000 1061.590 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.110 0.000 1075.390 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.370 0.000 1089.650 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.170 0.000 1103.450 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.970 0.000 1117.250 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.230 0.000 1131.510 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.030 0.000 1145.310 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 0.000 1159.570 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.090 0.000 1173.370 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.350 0.000 1187.630 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 0.000 1201.430 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.950 0.000 1215.230 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.210 0.000 1229.490 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.010 0.000 1243.290 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.270 0.000 1257.550 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.070 0.000 1271.350 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.330 0.000 1285.610 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.130 0.000 1299.410 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.930 0.000 1313.210 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.190 0.000 1327.470 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.990 0.000 1341.270 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.250 0.000 1355.530 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.050 0.000 1369.330 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1383.310 0.000 1383.590 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.110 0.000 1397.390 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.910 0.000 1411.190 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1425.170 0.000 1425.450 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.970 0.000 1439.250 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.230 0.000 1453.510 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.030 0.000 1467.310 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.290 0.000 1481.570 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.090 0.000 1495.370 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.890 0.000 1509.170 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.150 0.000 1523.430 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.950 0.000 1537.230 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.210 0.000 1551.490 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.010 0.000 1565.290 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.810 0.000 1579.090 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.070 0.000 1593.350 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.870 0.000 1607.150 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.130 0.000 1621.410 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.930 0.000 1635.210 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1649.190 0.000 1649.470 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.990 0.000 1663.270 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1676.790 0.000 1677.070 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.050 0.000 1691.330 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.850 0.000 1705.130 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.110 0.000 1719.390 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.910 0.000 1733.190 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.170 0.000 1747.450 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 0.000 613.550 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.970 0.000 1761.250 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.770 0.000 1775.050 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1789.030 0.000 1789.310 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1802.830 0.000 1803.110 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.090 0.000 1817.370 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1830.890 0.000 1831.170 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.150 0.000 1845.430 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.950 0.000 1859.230 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1872.750 0.000 1873.030 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.010 0.000 1887.290 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.410 0.000 1905.690 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1919.670 0.000 1919.950 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.470 0.000 1933.750 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.730 0.000 1948.010 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.530 0.000 1961.810 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1975.790 0.000 1976.070 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1989.590 0.000 1989.870 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.390 0.000 2003.670 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.650 0.000 2017.930 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2031.450 0.000 2031.730 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2045.710 0.000 2045.990 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.510 0.000 2059.790 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2073.770 0.000 2074.050 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2087.570 0.000 2087.850 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2101.370 0.000 2101.650 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2115.630 0.000 2115.910 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2129.430 0.000 2129.710 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2143.690 0.000 2143.970 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2157.490 0.000 2157.770 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2171.750 0.000 2172.030 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2185.550 0.000 2185.830 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2199.350 0.000 2199.630 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.610 0.000 2213.890 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2227.410 0.000 2227.690 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2241.670 0.000 2241.950 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2255.470 0.000 2255.750 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2269.730 0.000 2270.010 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2283.530 0.000 2283.810 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 0.000 674.270 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.790 0.000 688.070 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 0.000 702.330 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 0.000 716.130 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 0.000 730.390 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 0.000 758.450 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 0.000 772.250 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 0.000 520.170 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.030 0.000 800.310 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.830 0.000 814.110 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 0.000 828.370 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 0.000 842.170 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 0.000 855.970 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.950 0.000 870.230 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.750 0.000 884.030 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.010 0.000 898.290 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.810 0.000 912.090 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 0.000 534.430 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.070 0.000 926.350 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.870 0.000 940.150 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.670 0.000 953.950 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.930 0.000 968.210 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.730 0.000 982.010 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.990 0.000 996.270 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.790 0.000 1010.070 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 0.000 1024.330 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.850 0.000 1038.130 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.650 0.000 1051.930 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 0.000 548.230 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.910 0.000 1066.190 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.710 0.000 1079.990 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.970 0.000 1094.250 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 0.000 1108.050 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.030 0.000 1122.310 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1135.830 0.000 1136.110 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 0.000 1149.910 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.890 0.000 1164.170 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.690 0.000 1177.970 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.950 0.000 1192.230 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 0.000 562.490 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.750 0.000 1206.030 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.010 0.000 1220.290 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.810 0.000 1234.090 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.610 0.000 1247.890 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.870 0.000 1262.150 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.670 0.000 1275.950 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.930 0.000 1290.210 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.730 0.000 1304.010 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.990 0.000 1318.270 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1331.790 0.000 1332.070 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 0.000 576.290 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.590 0.000 1345.870 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.850 0.000 1360.130 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.650 0.000 1373.930 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.910 0.000 1388.190 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.710 0.000 1401.990 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.970 0.000 1416.250 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 0.000 1430.050 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.570 0.000 1443.850 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1457.830 0.000 1458.110 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 0.000 1471.910 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.890 0.000 1486.170 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.690 0.000 1499.970 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.950 0.000 1514.230 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.750 0.000 1528.030 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1541.550 0.000 1541.830 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.810 0.000 1556.090 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.610 0.000 1569.890 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.870 0.000 1584.150 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.670 0.000 1597.950 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.470 0.000 1611.750 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 0.000 604.350 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.730 0.000 1626.010 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.530 0.000 1639.810 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1653.790 0.000 1654.070 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.590 0.000 1667.870 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.850 0.000 1682.130 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1695.650 0.000 1695.930 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.450 0.000 1709.730 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1723.710 0.000 1723.990 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1737.510 0.000 1737.790 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.770 0.000 1752.050 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 0.000 618.150 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.570 0.000 1765.850 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1779.830 0.000 1780.110 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.630 0.000 1793.910 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1807.430 0.000 1807.710 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1821.690 0.000 1821.970 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.490 0.000 1835.770 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1849.750 0.000 1850.030 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1863.550 0.000 1863.830 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.810 0.000 1878.090 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1891.610 0.000 1891.890 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 0.000 632.410 4.000 ;
    END
  END la_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.040 10.640 122.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.040 10.640 522.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 721.040 10.640 722.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 821.040 10.640 822.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 10.640 922.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.040 10.640 1022.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.040 10.640 1122.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1221.040 10.640 1222.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1321.040 10.640 1322.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1421.040 10.640 1422.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1521.040 10.640 1522.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1621.040 10.640 1622.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.040 10.640 1722.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1821.040 10.640 1822.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1921.040 10.640 1922.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2021.040 10.640 2022.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2121.040 10.640 2122.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2221.040 10.640 2222.640 987.600 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 10.640 272.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.040 10.640 572.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.040 10.640 672.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 871.040 10.640 872.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 971.040 10.640 972.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 10.640 1072.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1171.040 10.640 1172.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1271.040 10.640 1272.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.040 10.640 1372.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1471.040 10.640 1472.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.040 10.640 1572.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1671.040 10.640 1672.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1771.040 10.640 1772.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1871.040 10.640 1872.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1971.040 10.640 1972.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2071.040 10.640 2072.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.040 10.640 2172.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2271.040 10.640 2272.640 987.600 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 0.000 343.070 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 0.000 441.050 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 0.000 454.850 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 0.000 482.910 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 0.000 277.750 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 0.000 361.470 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 0.000 445.650 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 0.000 487.510 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 0.000 464.510 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 0.000 478.310 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 0.000 492.110 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2294.480 987.445 ;
      LAYER met1 ;
        RECT 2.370 6.840 2297.630 987.600 ;
      LAYER met2 ;
        RECT 2.400 995.720 42.130 996.610 ;
        RECT 42.970 995.720 127.230 996.610 ;
        RECT 128.070 995.720 212.330 996.610 ;
        RECT 213.170 995.720 297.430 996.610 ;
        RECT 298.270 995.720 382.530 996.610 ;
        RECT 383.370 995.720 467.630 996.610 ;
        RECT 468.470 995.720 553.190 996.610 ;
        RECT 554.030 995.720 638.290 996.610 ;
        RECT 639.130 995.720 723.390 996.610 ;
        RECT 724.230 995.720 808.490 996.610 ;
        RECT 809.330 995.720 893.590 996.610 ;
        RECT 894.430 995.720 979.150 996.610 ;
        RECT 979.990 995.720 1064.250 996.610 ;
        RECT 1065.090 995.720 1149.350 996.610 ;
        RECT 1150.190 995.720 1234.450 996.610 ;
        RECT 1235.290 995.720 1319.550 996.610 ;
        RECT 1320.390 995.720 1404.650 996.610 ;
        RECT 1405.490 995.720 1490.210 996.610 ;
        RECT 1491.050 995.720 1575.310 996.610 ;
        RECT 1576.150 995.720 1660.410 996.610 ;
        RECT 1661.250 995.720 1745.510 996.610 ;
        RECT 1746.350 995.720 1830.610 996.610 ;
        RECT 1831.450 995.720 1916.170 996.610 ;
        RECT 1917.010 995.720 2001.270 996.610 ;
        RECT 2002.110 995.720 2086.370 996.610 ;
        RECT 2087.210 995.720 2171.470 996.610 ;
        RECT 2172.310 995.720 2256.570 996.610 ;
        RECT 2257.410 995.720 2297.600 996.610 ;
        RECT 2.400 4.280 2297.600 995.720 ;
        RECT 2.950 3.670 6.710 4.280 ;
        RECT 7.550 3.670 11.310 4.280 ;
        RECT 12.150 3.670 15.910 4.280 ;
        RECT 16.750 3.670 20.510 4.280 ;
        RECT 21.350 3.670 25.110 4.280 ;
        RECT 25.950 3.670 29.710 4.280 ;
        RECT 30.550 3.670 34.310 4.280 ;
        RECT 35.150 3.670 39.370 4.280 ;
        RECT 40.210 3.670 43.970 4.280 ;
        RECT 44.810 3.670 48.570 4.280 ;
        RECT 49.410 3.670 53.170 4.280 ;
        RECT 54.010 3.670 57.770 4.280 ;
        RECT 58.610 3.670 62.370 4.280 ;
        RECT 63.210 3.670 66.970 4.280 ;
        RECT 67.810 3.670 72.030 4.280 ;
        RECT 72.870 3.670 76.630 4.280 ;
        RECT 77.470 3.670 81.230 4.280 ;
        RECT 82.070 3.670 85.830 4.280 ;
        RECT 86.670 3.670 90.430 4.280 ;
        RECT 91.270 3.670 95.030 4.280 ;
        RECT 95.870 3.670 99.630 4.280 ;
        RECT 100.470 3.670 104.690 4.280 ;
        RECT 105.530 3.670 109.290 4.280 ;
        RECT 110.130 3.670 113.890 4.280 ;
        RECT 114.730 3.670 118.490 4.280 ;
        RECT 119.330 3.670 123.090 4.280 ;
        RECT 123.930 3.670 127.690 4.280 ;
        RECT 128.530 3.670 132.290 4.280 ;
        RECT 133.130 3.670 137.350 4.280 ;
        RECT 138.190 3.670 141.950 4.280 ;
        RECT 142.790 3.670 146.550 4.280 ;
        RECT 147.390 3.670 151.150 4.280 ;
        RECT 151.990 3.670 155.750 4.280 ;
        RECT 156.590 3.670 160.350 4.280 ;
        RECT 161.190 3.670 164.950 4.280 ;
        RECT 165.790 3.670 170.010 4.280 ;
        RECT 170.850 3.670 174.610 4.280 ;
        RECT 175.450 3.670 179.210 4.280 ;
        RECT 180.050 3.670 183.810 4.280 ;
        RECT 184.650 3.670 188.410 4.280 ;
        RECT 189.250 3.670 193.010 4.280 ;
        RECT 193.850 3.670 197.610 4.280 ;
        RECT 198.450 3.670 202.670 4.280 ;
        RECT 203.510 3.670 207.270 4.280 ;
        RECT 208.110 3.670 211.870 4.280 ;
        RECT 212.710 3.670 216.470 4.280 ;
        RECT 217.310 3.670 221.070 4.280 ;
        RECT 221.910 3.670 225.670 4.280 ;
        RECT 226.510 3.670 230.270 4.280 ;
        RECT 231.110 3.670 235.330 4.280 ;
        RECT 236.170 3.670 239.930 4.280 ;
        RECT 240.770 3.670 244.530 4.280 ;
        RECT 245.370 3.670 249.130 4.280 ;
        RECT 249.970 3.670 253.730 4.280 ;
        RECT 254.570 3.670 258.330 4.280 ;
        RECT 259.170 3.670 262.930 4.280 ;
        RECT 263.770 3.670 267.990 4.280 ;
        RECT 268.830 3.670 272.590 4.280 ;
        RECT 273.430 3.670 277.190 4.280 ;
        RECT 278.030 3.670 281.790 4.280 ;
        RECT 282.630 3.670 286.390 4.280 ;
        RECT 287.230 3.670 290.990 4.280 ;
        RECT 291.830 3.670 295.590 4.280 ;
        RECT 296.430 3.670 300.650 4.280 ;
        RECT 301.490 3.670 305.250 4.280 ;
        RECT 306.090 3.670 309.850 4.280 ;
        RECT 310.690 3.670 314.450 4.280 ;
        RECT 315.290 3.670 319.050 4.280 ;
        RECT 319.890 3.670 323.650 4.280 ;
        RECT 324.490 3.670 328.250 4.280 ;
        RECT 329.090 3.670 333.310 4.280 ;
        RECT 334.150 3.670 337.910 4.280 ;
        RECT 338.750 3.670 342.510 4.280 ;
        RECT 343.350 3.670 347.110 4.280 ;
        RECT 347.950 3.670 351.710 4.280 ;
        RECT 352.550 3.670 356.310 4.280 ;
        RECT 357.150 3.670 360.910 4.280 ;
        RECT 361.750 3.670 365.970 4.280 ;
        RECT 366.810 3.670 370.570 4.280 ;
        RECT 371.410 3.670 375.170 4.280 ;
        RECT 376.010 3.670 379.770 4.280 ;
        RECT 380.610 3.670 384.370 4.280 ;
        RECT 385.210 3.670 388.970 4.280 ;
        RECT 389.810 3.670 393.570 4.280 ;
        RECT 394.410 3.670 398.630 4.280 ;
        RECT 399.470 3.670 403.230 4.280 ;
        RECT 404.070 3.670 407.830 4.280 ;
        RECT 408.670 3.670 412.430 4.280 ;
        RECT 413.270 3.670 417.030 4.280 ;
        RECT 417.870 3.670 421.630 4.280 ;
        RECT 422.470 3.670 426.230 4.280 ;
        RECT 427.070 3.670 431.290 4.280 ;
        RECT 432.130 3.670 435.890 4.280 ;
        RECT 436.730 3.670 440.490 4.280 ;
        RECT 441.330 3.670 445.090 4.280 ;
        RECT 445.930 3.670 449.690 4.280 ;
        RECT 450.530 3.670 454.290 4.280 ;
        RECT 455.130 3.670 458.890 4.280 ;
        RECT 459.730 3.670 463.950 4.280 ;
        RECT 464.790 3.670 468.550 4.280 ;
        RECT 469.390 3.670 473.150 4.280 ;
        RECT 473.990 3.670 477.750 4.280 ;
        RECT 478.590 3.670 482.350 4.280 ;
        RECT 483.190 3.670 486.950 4.280 ;
        RECT 487.790 3.670 491.550 4.280 ;
        RECT 492.390 3.670 496.610 4.280 ;
        RECT 497.450 3.670 501.210 4.280 ;
        RECT 502.050 3.670 505.810 4.280 ;
        RECT 506.650 3.670 510.410 4.280 ;
        RECT 511.250 3.670 515.010 4.280 ;
        RECT 515.850 3.670 519.610 4.280 ;
        RECT 520.450 3.670 524.210 4.280 ;
        RECT 525.050 3.670 529.270 4.280 ;
        RECT 530.110 3.670 533.870 4.280 ;
        RECT 534.710 3.670 538.470 4.280 ;
        RECT 539.310 3.670 543.070 4.280 ;
        RECT 543.910 3.670 547.670 4.280 ;
        RECT 548.510 3.670 552.270 4.280 ;
        RECT 553.110 3.670 556.870 4.280 ;
        RECT 557.710 3.670 561.930 4.280 ;
        RECT 562.770 3.670 566.530 4.280 ;
        RECT 567.370 3.670 571.130 4.280 ;
        RECT 571.970 3.670 575.730 4.280 ;
        RECT 576.570 3.670 580.330 4.280 ;
        RECT 581.170 3.670 584.930 4.280 ;
        RECT 585.770 3.670 589.530 4.280 ;
        RECT 590.370 3.670 594.590 4.280 ;
        RECT 595.430 3.670 599.190 4.280 ;
        RECT 600.030 3.670 603.790 4.280 ;
        RECT 604.630 3.670 608.390 4.280 ;
        RECT 609.230 3.670 612.990 4.280 ;
        RECT 613.830 3.670 617.590 4.280 ;
        RECT 618.430 3.670 622.190 4.280 ;
        RECT 623.030 3.670 627.250 4.280 ;
        RECT 628.090 3.670 631.850 4.280 ;
        RECT 632.690 3.670 636.450 4.280 ;
        RECT 637.290 3.670 641.050 4.280 ;
        RECT 641.890 3.670 645.650 4.280 ;
        RECT 646.490 3.670 650.250 4.280 ;
        RECT 651.090 3.670 654.850 4.280 ;
        RECT 655.690 3.670 659.910 4.280 ;
        RECT 660.750 3.670 664.510 4.280 ;
        RECT 665.350 3.670 669.110 4.280 ;
        RECT 669.950 3.670 673.710 4.280 ;
        RECT 674.550 3.670 678.310 4.280 ;
        RECT 679.150 3.670 682.910 4.280 ;
        RECT 683.750 3.670 687.510 4.280 ;
        RECT 688.350 3.670 692.570 4.280 ;
        RECT 693.410 3.670 697.170 4.280 ;
        RECT 698.010 3.670 701.770 4.280 ;
        RECT 702.610 3.670 706.370 4.280 ;
        RECT 707.210 3.670 710.970 4.280 ;
        RECT 711.810 3.670 715.570 4.280 ;
        RECT 716.410 3.670 720.170 4.280 ;
        RECT 721.010 3.670 725.230 4.280 ;
        RECT 726.070 3.670 729.830 4.280 ;
        RECT 730.670 3.670 734.430 4.280 ;
        RECT 735.270 3.670 739.030 4.280 ;
        RECT 739.870 3.670 743.630 4.280 ;
        RECT 744.470 3.670 748.230 4.280 ;
        RECT 749.070 3.670 752.830 4.280 ;
        RECT 753.670 3.670 757.890 4.280 ;
        RECT 758.730 3.670 762.490 4.280 ;
        RECT 763.330 3.670 767.090 4.280 ;
        RECT 767.930 3.670 771.690 4.280 ;
        RECT 772.530 3.670 776.290 4.280 ;
        RECT 777.130 3.670 780.890 4.280 ;
        RECT 781.730 3.670 785.490 4.280 ;
        RECT 786.330 3.670 790.090 4.280 ;
        RECT 790.930 3.670 795.150 4.280 ;
        RECT 795.990 3.670 799.750 4.280 ;
        RECT 800.590 3.670 804.350 4.280 ;
        RECT 805.190 3.670 808.950 4.280 ;
        RECT 809.790 3.670 813.550 4.280 ;
        RECT 814.390 3.670 818.150 4.280 ;
        RECT 818.990 3.670 822.750 4.280 ;
        RECT 823.590 3.670 827.810 4.280 ;
        RECT 828.650 3.670 832.410 4.280 ;
        RECT 833.250 3.670 837.010 4.280 ;
        RECT 837.850 3.670 841.610 4.280 ;
        RECT 842.450 3.670 846.210 4.280 ;
        RECT 847.050 3.670 850.810 4.280 ;
        RECT 851.650 3.670 855.410 4.280 ;
        RECT 856.250 3.670 860.470 4.280 ;
        RECT 861.310 3.670 865.070 4.280 ;
        RECT 865.910 3.670 869.670 4.280 ;
        RECT 870.510 3.670 874.270 4.280 ;
        RECT 875.110 3.670 878.870 4.280 ;
        RECT 879.710 3.670 883.470 4.280 ;
        RECT 884.310 3.670 888.070 4.280 ;
        RECT 888.910 3.670 893.130 4.280 ;
        RECT 893.970 3.670 897.730 4.280 ;
        RECT 898.570 3.670 902.330 4.280 ;
        RECT 903.170 3.670 906.930 4.280 ;
        RECT 907.770 3.670 911.530 4.280 ;
        RECT 912.370 3.670 916.130 4.280 ;
        RECT 916.970 3.670 920.730 4.280 ;
        RECT 921.570 3.670 925.790 4.280 ;
        RECT 926.630 3.670 930.390 4.280 ;
        RECT 931.230 3.670 934.990 4.280 ;
        RECT 935.830 3.670 939.590 4.280 ;
        RECT 940.430 3.670 944.190 4.280 ;
        RECT 945.030 3.670 948.790 4.280 ;
        RECT 949.630 3.670 953.390 4.280 ;
        RECT 954.230 3.670 958.450 4.280 ;
        RECT 959.290 3.670 963.050 4.280 ;
        RECT 963.890 3.670 967.650 4.280 ;
        RECT 968.490 3.670 972.250 4.280 ;
        RECT 973.090 3.670 976.850 4.280 ;
        RECT 977.690 3.670 981.450 4.280 ;
        RECT 982.290 3.670 986.050 4.280 ;
        RECT 986.890 3.670 991.110 4.280 ;
        RECT 991.950 3.670 995.710 4.280 ;
        RECT 996.550 3.670 1000.310 4.280 ;
        RECT 1001.150 3.670 1004.910 4.280 ;
        RECT 1005.750 3.670 1009.510 4.280 ;
        RECT 1010.350 3.670 1014.110 4.280 ;
        RECT 1014.950 3.670 1018.710 4.280 ;
        RECT 1019.550 3.670 1023.770 4.280 ;
        RECT 1024.610 3.670 1028.370 4.280 ;
        RECT 1029.210 3.670 1032.970 4.280 ;
        RECT 1033.810 3.670 1037.570 4.280 ;
        RECT 1038.410 3.670 1042.170 4.280 ;
        RECT 1043.010 3.670 1046.770 4.280 ;
        RECT 1047.610 3.670 1051.370 4.280 ;
        RECT 1052.210 3.670 1056.430 4.280 ;
        RECT 1057.270 3.670 1061.030 4.280 ;
        RECT 1061.870 3.670 1065.630 4.280 ;
        RECT 1066.470 3.670 1070.230 4.280 ;
        RECT 1071.070 3.670 1074.830 4.280 ;
        RECT 1075.670 3.670 1079.430 4.280 ;
        RECT 1080.270 3.670 1084.030 4.280 ;
        RECT 1084.870 3.670 1089.090 4.280 ;
        RECT 1089.930 3.670 1093.690 4.280 ;
        RECT 1094.530 3.670 1098.290 4.280 ;
        RECT 1099.130 3.670 1102.890 4.280 ;
        RECT 1103.730 3.670 1107.490 4.280 ;
        RECT 1108.330 3.670 1112.090 4.280 ;
        RECT 1112.930 3.670 1116.690 4.280 ;
        RECT 1117.530 3.670 1121.750 4.280 ;
        RECT 1122.590 3.670 1126.350 4.280 ;
        RECT 1127.190 3.670 1130.950 4.280 ;
        RECT 1131.790 3.670 1135.550 4.280 ;
        RECT 1136.390 3.670 1140.150 4.280 ;
        RECT 1140.990 3.670 1144.750 4.280 ;
        RECT 1145.590 3.670 1149.350 4.280 ;
        RECT 1150.190 3.670 1154.410 4.280 ;
        RECT 1155.250 3.670 1159.010 4.280 ;
        RECT 1159.850 3.670 1163.610 4.280 ;
        RECT 1164.450 3.670 1168.210 4.280 ;
        RECT 1169.050 3.670 1172.810 4.280 ;
        RECT 1173.650 3.670 1177.410 4.280 ;
        RECT 1178.250 3.670 1182.010 4.280 ;
        RECT 1182.850 3.670 1187.070 4.280 ;
        RECT 1187.910 3.670 1191.670 4.280 ;
        RECT 1192.510 3.670 1196.270 4.280 ;
        RECT 1197.110 3.670 1200.870 4.280 ;
        RECT 1201.710 3.670 1205.470 4.280 ;
        RECT 1206.310 3.670 1210.070 4.280 ;
        RECT 1210.910 3.670 1214.670 4.280 ;
        RECT 1215.510 3.670 1219.730 4.280 ;
        RECT 1220.570 3.670 1224.330 4.280 ;
        RECT 1225.170 3.670 1228.930 4.280 ;
        RECT 1229.770 3.670 1233.530 4.280 ;
        RECT 1234.370 3.670 1238.130 4.280 ;
        RECT 1238.970 3.670 1242.730 4.280 ;
        RECT 1243.570 3.670 1247.330 4.280 ;
        RECT 1248.170 3.670 1252.390 4.280 ;
        RECT 1253.230 3.670 1256.990 4.280 ;
        RECT 1257.830 3.670 1261.590 4.280 ;
        RECT 1262.430 3.670 1266.190 4.280 ;
        RECT 1267.030 3.670 1270.790 4.280 ;
        RECT 1271.630 3.670 1275.390 4.280 ;
        RECT 1276.230 3.670 1279.990 4.280 ;
        RECT 1280.830 3.670 1285.050 4.280 ;
        RECT 1285.890 3.670 1289.650 4.280 ;
        RECT 1290.490 3.670 1294.250 4.280 ;
        RECT 1295.090 3.670 1298.850 4.280 ;
        RECT 1299.690 3.670 1303.450 4.280 ;
        RECT 1304.290 3.670 1308.050 4.280 ;
        RECT 1308.890 3.670 1312.650 4.280 ;
        RECT 1313.490 3.670 1317.710 4.280 ;
        RECT 1318.550 3.670 1322.310 4.280 ;
        RECT 1323.150 3.670 1326.910 4.280 ;
        RECT 1327.750 3.670 1331.510 4.280 ;
        RECT 1332.350 3.670 1336.110 4.280 ;
        RECT 1336.950 3.670 1340.710 4.280 ;
        RECT 1341.550 3.670 1345.310 4.280 ;
        RECT 1346.150 3.670 1350.370 4.280 ;
        RECT 1351.210 3.670 1354.970 4.280 ;
        RECT 1355.810 3.670 1359.570 4.280 ;
        RECT 1360.410 3.670 1364.170 4.280 ;
        RECT 1365.010 3.670 1368.770 4.280 ;
        RECT 1369.610 3.670 1373.370 4.280 ;
        RECT 1374.210 3.670 1377.970 4.280 ;
        RECT 1378.810 3.670 1383.030 4.280 ;
        RECT 1383.870 3.670 1387.630 4.280 ;
        RECT 1388.470 3.670 1392.230 4.280 ;
        RECT 1393.070 3.670 1396.830 4.280 ;
        RECT 1397.670 3.670 1401.430 4.280 ;
        RECT 1402.270 3.670 1406.030 4.280 ;
        RECT 1406.870 3.670 1410.630 4.280 ;
        RECT 1411.470 3.670 1415.690 4.280 ;
        RECT 1416.530 3.670 1420.290 4.280 ;
        RECT 1421.130 3.670 1424.890 4.280 ;
        RECT 1425.730 3.670 1429.490 4.280 ;
        RECT 1430.330 3.670 1434.090 4.280 ;
        RECT 1434.930 3.670 1438.690 4.280 ;
        RECT 1439.530 3.670 1443.290 4.280 ;
        RECT 1444.130 3.670 1448.350 4.280 ;
        RECT 1449.190 3.670 1452.950 4.280 ;
        RECT 1453.790 3.670 1457.550 4.280 ;
        RECT 1458.390 3.670 1462.150 4.280 ;
        RECT 1462.990 3.670 1466.750 4.280 ;
        RECT 1467.590 3.670 1471.350 4.280 ;
        RECT 1472.190 3.670 1475.950 4.280 ;
        RECT 1476.790 3.670 1481.010 4.280 ;
        RECT 1481.850 3.670 1485.610 4.280 ;
        RECT 1486.450 3.670 1490.210 4.280 ;
        RECT 1491.050 3.670 1494.810 4.280 ;
        RECT 1495.650 3.670 1499.410 4.280 ;
        RECT 1500.250 3.670 1504.010 4.280 ;
        RECT 1504.850 3.670 1508.610 4.280 ;
        RECT 1509.450 3.670 1513.670 4.280 ;
        RECT 1514.510 3.670 1518.270 4.280 ;
        RECT 1519.110 3.670 1522.870 4.280 ;
        RECT 1523.710 3.670 1527.470 4.280 ;
        RECT 1528.310 3.670 1532.070 4.280 ;
        RECT 1532.910 3.670 1536.670 4.280 ;
        RECT 1537.510 3.670 1541.270 4.280 ;
        RECT 1542.110 3.670 1545.870 4.280 ;
        RECT 1546.710 3.670 1550.930 4.280 ;
        RECT 1551.770 3.670 1555.530 4.280 ;
        RECT 1556.370 3.670 1560.130 4.280 ;
        RECT 1560.970 3.670 1564.730 4.280 ;
        RECT 1565.570 3.670 1569.330 4.280 ;
        RECT 1570.170 3.670 1573.930 4.280 ;
        RECT 1574.770 3.670 1578.530 4.280 ;
        RECT 1579.370 3.670 1583.590 4.280 ;
        RECT 1584.430 3.670 1588.190 4.280 ;
        RECT 1589.030 3.670 1592.790 4.280 ;
        RECT 1593.630 3.670 1597.390 4.280 ;
        RECT 1598.230 3.670 1601.990 4.280 ;
        RECT 1602.830 3.670 1606.590 4.280 ;
        RECT 1607.430 3.670 1611.190 4.280 ;
        RECT 1612.030 3.670 1616.250 4.280 ;
        RECT 1617.090 3.670 1620.850 4.280 ;
        RECT 1621.690 3.670 1625.450 4.280 ;
        RECT 1626.290 3.670 1630.050 4.280 ;
        RECT 1630.890 3.670 1634.650 4.280 ;
        RECT 1635.490 3.670 1639.250 4.280 ;
        RECT 1640.090 3.670 1643.850 4.280 ;
        RECT 1644.690 3.670 1648.910 4.280 ;
        RECT 1649.750 3.670 1653.510 4.280 ;
        RECT 1654.350 3.670 1658.110 4.280 ;
        RECT 1658.950 3.670 1662.710 4.280 ;
        RECT 1663.550 3.670 1667.310 4.280 ;
        RECT 1668.150 3.670 1671.910 4.280 ;
        RECT 1672.750 3.670 1676.510 4.280 ;
        RECT 1677.350 3.670 1681.570 4.280 ;
        RECT 1682.410 3.670 1686.170 4.280 ;
        RECT 1687.010 3.670 1690.770 4.280 ;
        RECT 1691.610 3.670 1695.370 4.280 ;
        RECT 1696.210 3.670 1699.970 4.280 ;
        RECT 1700.810 3.670 1704.570 4.280 ;
        RECT 1705.410 3.670 1709.170 4.280 ;
        RECT 1710.010 3.670 1714.230 4.280 ;
        RECT 1715.070 3.670 1718.830 4.280 ;
        RECT 1719.670 3.670 1723.430 4.280 ;
        RECT 1724.270 3.670 1728.030 4.280 ;
        RECT 1728.870 3.670 1732.630 4.280 ;
        RECT 1733.470 3.670 1737.230 4.280 ;
        RECT 1738.070 3.670 1741.830 4.280 ;
        RECT 1742.670 3.670 1746.890 4.280 ;
        RECT 1747.730 3.670 1751.490 4.280 ;
        RECT 1752.330 3.670 1756.090 4.280 ;
        RECT 1756.930 3.670 1760.690 4.280 ;
        RECT 1761.530 3.670 1765.290 4.280 ;
        RECT 1766.130 3.670 1769.890 4.280 ;
        RECT 1770.730 3.670 1774.490 4.280 ;
        RECT 1775.330 3.670 1779.550 4.280 ;
        RECT 1780.390 3.670 1784.150 4.280 ;
        RECT 1784.990 3.670 1788.750 4.280 ;
        RECT 1789.590 3.670 1793.350 4.280 ;
        RECT 1794.190 3.670 1797.950 4.280 ;
        RECT 1798.790 3.670 1802.550 4.280 ;
        RECT 1803.390 3.670 1807.150 4.280 ;
        RECT 1807.990 3.670 1812.210 4.280 ;
        RECT 1813.050 3.670 1816.810 4.280 ;
        RECT 1817.650 3.670 1821.410 4.280 ;
        RECT 1822.250 3.670 1826.010 4.280 ;
        RECT 1826.850 3.670 1830.610 4.280 ;
        RECT 1831.450 3.670 1835.210 4.280 ;
        RECT 1836.050 3.670 1839.810 4.280 ;
        RECT 1840.650 3.670 1844.870 4.280 ;
        RECT 1845.710 3.670 1849.470 4.280 ;
        RECT 1850.310 3.670 1854.070 4.280 ;
        RECT 1854.910 3.670 1858.670 4.280 ;
        RECT 1859.510 3.670 1863.270 4.280 ;
        RECT 1864.110 3.670 1867.870 4.280 ;
        RECT 1868.710 3.670 1872.470 4.280 ;
        RECT 1873.310 3.670 1877.530 4.280 ;
        RECT 1878.370 3.670 1882.130 4.280 ;
        RECT 1882.970 3.670 1886.730 4.280 ;
        RECT 1887.570 3.670 1891.330 4.280 ;
        RECT 1892.170 3.670 1895.930 4.280 ;
        RECT 1896.770 3.670 1900.530 4.280 ;
        RECT 1901.370 3.670 1905.130 4.280 ;
        RECT 1905.970 3.670 1910.190 4.280 ;
        RECT 1911.030 3.670 1914.790 4.280 ;
        RECT 1915.630 3.670 1919.390 4.280 ;
        RECT 1920.230 3.670 1923.990 4.280 ;
        RECT 1924.830 3.670 1928.590 4.280 ;
        RECT 1929.430 3.670 1933.190 4.280 ;
        RECT 1934.030 3.670 1937.790 4.280 ;
        RECT 1938.630 3.670 1942.850 4.280 ;
        RECT 1943.690 3.670 1947.450 4.280 ;
        RECT 1948.290 3.670 1952.050 4.280 ;
        RECT 1952.890 3.670 1956.650 4.280 ;
        RECT 1957.490 3.670 1961.250 4.280 ;
        RECT 1962.090 3.670 1965.850 4.280 ;
        RECT 1966.690 3.670 1970.450 4.280 ;
        RECT 1971.290 3.670 1975.510 4.280 ;
        RECT 1976.350 3.670 1980.110 4.280 ;
        RECT 1980.950 3.670 1984.710 4.280 ;
        RECT 1985.550 3.670 1989.310 4.280 ;
        RECT 1990.150 3.670 1993.910 4.280 ;
        RECT 1994.750 3.670 1998.510 4.280 ;
        RECT 1999.350 3.670 2003.110 4.280 ;
        RECT 2003.950 3.670 2008.170 4.280 ;
        RECT 2009.010 3.670 2012.770 4.280 ;
        RECT 2013.610 3.670 2017.370 4.280 ;
        RECT 2018.210 3.670 2021.970 4.280 ;
        RECT 2022.810 3.670 2026.570 4.280 ;
        RECT 2027.410 3.670 2031.170 4.280 ;
        RECT 2032.010 3.670 2035.770 4.280 ;
        RECT 2036.610 3.670 2040.830 4.280 ;
        RECT 2041.670 3.670 2045.430 4.280 ;
        RECT 2046.270 3.670 2050.030 4.280 ;
        RECT 2050.870 3.670 2054.630 4.280 ;
        RECT 2055.470 3.670 2059.230 4.280 ;
        RECT 2060.070 3.670 2063.830 4.280 ;
        RECT 2064.670 3.670 2068.430 4.280 ;
        RECT 2069.270 3.670 2073.490 4.280 ;
        RECT 2074.330 3.670 2078.090 4.280 ;
        RECT 2078.930 3.670 2082.690 4.280 ;
        RECT 2083.530 3.670 2087.290 4.280 ;
        RECT 2088.130 3.670 2091.890 4.280 ;
        RECT 2092.730 3.670 2096.490 4.280 ;
        RECT 2097.330 3.670 2101.090 4.280 ;
        RECT 2101.930 3.670 2106.150 4.280 ;
        RECT 2106.990 3.670 2110.750 4.280 ;
        RECT 2111.590 3.670 2115.350 4.280 ;
        RECT 2116.190 3.670 2119.950 4.280 ;
        RECT 2120.790 3.670 2124.550 4.280 ;
        RECT 2125.390 3.670 2129.150 4.280 ;
        RECT 2129.990 3.670 2133.750 4.280 ;
        RECT 2134.590 3.670 2138.810 4.280 ;
        RECT 2139.650 3.670 2143.410 4.280 ;
        RECT 2144.250 3.670 2148.010 4.280 ;
        RECT 2148.850 3.670 2152.610 4.280 ;
        RECT 2153.450 3.670 2157.210 4.280 ;
        RECT 2158.050 3.670 2161.810 4.280 ;
        RECT 2162.650 3.670 2166.410 4.280 ;
        RECT 2167.250 3.670 2171.470 4.280 ;
        RECT 2172.310 3.670 2176.070 4.280 ;
        RECT 2176.910 3.670 2180.670 4.280 ;
        RECT 2181.510 3.670 2185.270 4.280 ;
        RECT 2186.110 3.670 2189.870 4.280 ;
        RECT 2190.710 3.670 2194.470 4.280 ;
        RECT 2195.310 3.670 2199.070 4.280 ;
        RECT 2199.910 3.670 2204.130 4.280 ;
        RECT 2204.970 3.670 2208.730 4.280 ;
        RECT 2209.570 3.670 2213.330 4.280 ;
        RECT 2214.170 3.670 2217.930 4.280 ;
        RECT 2218.770 3.670 2222.530 4.280 ;
        RECT 2223.370 3.670 2227.130 4.280 ;
        RECT 2227.970 3.670 2231.730 4.280 ;
        RECT 2232.570 3.670 2236.790 4.280 ;
        RECT 2237.630 3.670 2241.390 4.280 ;
        RECT 2242.230 3.670 2245.990 4.280 ;
        RECT 2246.830 3.670 2250.590 4.280 ;
        RECT 2251.430 3.670 2255.190 4.280 ;
        RECT 2256.030 3.670 2259.790 4.280 ;
        RECT 2260.630 3.670 2264.390 4.280 ;
        RECT 2265.230 3.670 2269.450 4.280 ;
        RECT 2270.290 3.670 2274.050 4.280 ;
        RECT 2274.890 3.670 2278.650 4.280 ;
        RECT 2279.490 3.670 2283.250 4.280 ;
        RECT 2284.090 3.670 2287.850 4.280 ;
        RECT 2288.690 3.670 2292.450 4.280 ;
        RECT 2293.290 3.670 2297.050 4.280 ;
      LAYER met3 ;
        RECT 4.000 988.400 2295.600 989.225 ;
        RECT 4.400 988.360 2295.600 988.400 ;
        RECT 4.400 987.000 2296.000 988.360 ;
        RECT 4.000 967.320 2296.000 987.000 ;
        RECT 4.000 965.920 2295.600 967.320 ;
        RECT 4.000 964.600 2296.000 965.920 ;
        RECT 4.400 963.200 2296.000 964.600 ;
        RECT 4.000 944.880 2296.000 963.200 ;
        RECT 4.000 943.480 2295.600 944.880 ;
        RECT 4.000 940.800 2296.000 943.480 ;
        RECT 4.400 939.400 2296.000 940.800 ;
        RECT 4.000 923.120 2296.000 939.400 ;
        RECT 4.000 921.720 2295.600 923.120 ;
        RECT 4.000 917.000 2296.000 921.720 ;
        RECT 4.400 915.600 2296.000 917.000 ;
        RECT 4.000 900.680 2296.000 915.600 ;
        RECT 4.000 899.280 2295.600 900.680 ;
        RECT 4.000 893.200 2296.000 899.280 ;
        RECT 4.400 891.800 2296.000 893.200 ;
        RECT 4.000 878.240 2296.000 891.800 ;
        RECT 4.000 876.840 2295.600 878.240 ;
        RECT 4.000 869.400 2296.000 876.840 ;
        RECT 4.400 868.000 2296.000 869.400 ;
        RECT 4.000 856.480 2296.000 868.000 ;
        RECT 4.000 855.080 2295.600 856.480 ;
        RECT 4.000 845.600 2296.000 855.080 ;
        RECT 4.400 844.200 2296.000 845.600 ;
        RECT 4.000 834.040 2296.000 844.200 ;
        RECT 4.000 832.640 2295.600 834.040 ;
        RECT 4.000 821.800 2296.000 832.640 ;
        RECT 4.400 820.400 2296.000 821.800 ;
        RECT 4.000 811.600 2296.000 820.400 ;
        RECT 4.000 810.200 2295.600 811.600 ;
        RECT 4.000 798.000 2296.000 810.200 ;
        RECT 4.400 796.600 2296.000 798.000 ;
        RECT 4.000 789.840 2296.000 796.600 ;
        RECT 4.000 788.440 2295.600 789.840 ;
        RECT 4.000 774.200 2296.000 788.440 ;
        RECT 4.400 772.800 2296.000 774.200 ;
        RECT 4.000 767.400 2296.000 772.800 ;
        RECT 4.000 766.000 2295.600 767.400 ;
        RECT 4.000 750.400 2296.000 766.000 ;
        RECT 4.400 749.000 2296.000 750.400 ;
        RECT 4.000 744.960 2296.000 749.000 ;
        RECT 4.000 743.560 2295.600 744.960 ;
        RECT 4.000 726.600 2296.000 743.560 ;
        RECT 4.400 725.200 2296.000 726.600 ;
        RECT 4.000 723.200 2296.000 725.200 ;
        RECT 4.000 721.800 2295.600 723.200 ;
        RECT 4.000 702.800 2296.000 721.800 ;
        RECT 4.400 701.400 2296.000 702.800 ;
        RECT 4.000 700.760 2296.000 701.400 ;
        RECT 4.000 699.360 2295.600 700.760 ;
        RECT 4.000 679.000 2296.000 699.360 ;
        RECT 4.400 678.320 2296.000 679.000 ;
        RECT 4.400 677.600 2295.600 678.320 ;
        RECT 4.000 676.920 2295.600 677.600 ;
        RECT 4.000 655.880 2296.000 676.920 ;
        RECT 4.000 655.200 2295.600 655.880 ;
        RECT 4.400 654.480 2295.600 655.200 ;
        RECT 4.400 653.800 2296.000 654.480 ;
        RECT 4.000 634.120 2296.000 653.800 ;
        RECT 4.000 632.720 2295.600 634.120 ;
        RECT 4.000 631.400 2296.000 632.720 ;
        RECT 4.400 630.000 2296.000 631.400 ;
        RECT 4.000 611.680 2296.000 630.000 ;
        RECT 4.000 610.280 2295.600 611.680 ;
        RECT 4.000 607.600 2296.000 610.280 ;
        RECT 4.400 606.200 2296.000 607.600 ;
        RECT 4.000 589.240 2296.000 606.200 ;
        RECT 4.000 587.840 2295.600 589.240 ;
        RECT 4.000 583.800 2296.000 587.840 ;
        RECT 4.400 582.400 2296.000 583.800 ;
        RECT 4.000 567.480 2296.000 582.400 ;
        RECT 4.000 566.080 2295.600 567.480 ;
        RECT 4.000 560.000 2296.000 566.080 ;
        RECT 4.400 558.600 2296.000 560.000 ;
        RECT 4.000 545.040 2296.000 558.600 ;
        RECT 4.000 543.640 2295.600 545.040 ;
        RECT 4.000 536.200 2296.000 543.640 ;
        RECT 4.400 534.800 2296.000 536.200 ;
        RECT 4.000 522.600 2296.000 534.800 ;
        RECT 4.000 521.200 2295.600 522.600 ;
        RECT 4.000 512.400 2296.000 521.200 ;
        RECT 4.400 511.000 2296.000 512.400 ;
        RECT 4.000 500.840 2296.000 511.000 ;
        RECT 4.000 499.440 2295.600 500.840 ;
        RECT 4.000 488.600 2296.000 499.440 ;
        RECT 4.400 487.200 2296.000 488.600 ;
        RECT 4.000 478.400 2296.000 487.200 ;
        RECT 4.000 477.000 2295.600 478.400 ;
        RECT 4.000 464.800 2296.000 477.000 ;
        RECT 4.400 463.400 2296.000 464.800 ;
        RECT 4.000 455.960 2296.000 463.400 ;
        RECT 4.000 454.560 2295.600 455.960 ;
        RECT 4.000 441.000 2296.000 454.560 ;
        RECT 4.400 439.600 2296.000 441.000 ;
        RECT 4.000 434.200 2296.000 439.600 ;
        RECT 4.000 432.800 2295.600 434.200 ;
        RECT 4.000 417.200 2296.000 432.800 ;
        RECT 4.400 415.800 2296.000 417.200 ;
        RECT 4.000 411.760 2296.000 415.800 ;
        RECT 4.000 410.360 2295.600 411.760 ;
        RECT 4.000 393.400 2296.000 410.360 ;
        RECT 4.400 392.000 2296.000 393.400 ;
        RECT 4.000 389.320 2296.000 392.000 ;
        RECT 4.000 387.920 2295.600 389.320 ;
        RECT 4.000 369.600 2296.000 387.920 ;
        RECT 4.400 368.200 2296.000 369.600 ;
        RECT 4.000 367.560 2296.000 368.200 ;
        RECT 4.000 366.160 2295.600 367.560 ;
        RECT 4.000 345.800 2296.000 366.160 ;
        RECT 4.400 345.120 2296.000 345.800 ;
        RECT 4.400 344.400 2295.600 345.120 ;
        RECT 4.000 343.720 2295.600 344.400 ;
        RECT 4.000 322.680 2296.000 343.720 ;
        RECT 4.000 322.000 2295.600 322.680 ;
        RECT 4.400 321.280 2295.600 322.000 ;
        RECT 4.400 320.600 2296.000 321.280 ;
        RECT 4.000 300.240 2296.000 320.600 ;
        RECT 4.000 298.840 2295.600 300.240 ;
        RECT 4.000 298.200 2296.000 298.840 ;
        RECT 4.400 296.800 2296.000 298.200 ;
        RECT 4.000 278.480 2296.000 296.800 ;
        RECT 4.000 277.080 2295.600 278.480 ;
        RECT 4.000 274.400 2296.000 277.080 ;
        RECT 4.400 273.000 2296.000 274.400 ;
        RECT 4.000 256.040 2296.000 273.000 ;
        RECT 4.000 254.640 2295.600 256.040 ;
        RECT 4.000 250.600 2296.000 254.640 ;
        RECT 4.400 249.200 2296.000 250.600 ;
        RECT 4.000 233.600 2296.000 249.200 ;
        RECT 4.000 232.200 2295.600 233.600 ;
        RECT 4.000 226.800 2296.000 232.200 ;
        RECT 4.400 225.400 2296.000 226.800 ;
        RECT 4.000 211.840 2296.000 225.400 ;
        RECT 4.000 210.440 2295.600 211.840 ;
        RECT 4.000 203.000 2296.000 210.440 ;
        RECT 4.400 201.600 2296.000 203.000 ;
        RECT 4.000 189.400 2296.000 201.600 ;
        RECT 4.000 188.000 2295.600 189.400 ;
        RECT 4.000 179.200 2296.000 188.000 ;
        RECT 4.400 177.800 2296.000 179.200 ;
        RECT 4.000 166.960 2296.000 177.800 ;
        RECT 4.000 165.560 2295.600 166.960 ;
        RECT 4.000 155.400 2296.000 165.560 ;
        RECT 4.400 154.000 2296.000 155.400 ;
        RECT 4.000 145.200 2296.000 154.000 ;
        RECT 4.000 143.800 2295.600 145.200 ;
        RECT 4.000 131.600 2296.000 143.800 ;
        RECT 4.400 130.200 2296.000 131.600 ;
        RECT 4.000 122.760 2296.000 130.200 ;
        RECT 4.000 121.360 2295.600 122.760 ;
        RECT 4.000 107.800 2296.000 121.360 ;
        RECT 4.400 106.400 2296.000 107.800 ;
        RECT 4.000 100.320 2296.000 106.400 ;
        RECT 4.000 98.920 2295.600 100.320 ;
        RECT 4.000 84.000 2296.000 98.920 ;
        RECT 4.400 82.600 2296.000 84.000 ;
        RECT 4.000 78.560 2296.000 82.600 ;
        RECT 4.000 77.160 2295.600 78.560 ;
        RECT 4.000 60.200 2296.000 77.160 ;
        RECT 4.400 58.800 2296.000 60.200 ;
        RECT 4.000 56.120 2296.000 58.800 ;
        RECT 4.000 54.720 2295.600 56.120 ;
        RECT 4.000 36.400 2296.000 54.720 ;
        RECT 4.400 35.000 2296.000 36.400 ;
        RECT 4.000 33.680 2296.000 35.000 ;
        RECT 4.000 32.280 2295.600 33.680 ;
        RECT 4.000 12.600 2296.000 32.280 ;
        RECT 4.400 11.920 2296.000 12.600 ;
        RECT 4.400 11.200 2295.600 11.920 ;
        RECT 4.000 10.715 2295.600 11.200 ;
      LAYER met4 ;
        RECT 370.135 58.655 370.640 821.265 ;
        RECT 373.040 58.655 420.640 821.265 ;
        RECT 423.040 58.655 470.640 821.265 ;
        RECT 473.040 58.655 520.640 821.265 ;
        RECT 523.040 58.655 570.640 821.265 ;
        RECT 573.040 58.655 620.640 821.265 ;
        RECT 623.040 58.655 670.640 821.265 ;
        RECT 673.040 58.655 720.640 821.265 ;
        RECT 723.040 58.655 770.640 821.265 ;
        RECT 773.040 58.655 820.640 821.265 ;
        RECT 823.040 58.655 870.640 821.265 ;
        RECT 873.040 58.655 920.640 821.265 ;
        RECT 923.040 58.655 970.640 821.265 ;
        RECT 973.040 58.655 1020.640 821.265 ;
        RECT 1023.040 58.655 1070.640 821.265 ;
        RECT 1073.040 58.655 1120.640 821.265 ;
        RECT 1123.040 58.655 1170.640 821.265 ;
        RECT 1173.040 58.655 1220.640 821.265 ;
        RECT 1223.040 58.655 1270.640 821.265 ;
        RECT 1273.040 58.655 1320.640 821.265 ;
        RECT 1323.040 58.655 1370.640 821.265 ;
        RECT 1373.040 58.655 1420.640 821.265 ;
        RECT 1423.040 58.655 1470.640 821.265 ;
        RECT 1473.040 58.655 1520.640 821.265 ;
        RECT 1523.040 58.655 1570.640 821.265 ;
        RECT 1573.040 58.655 1620.640 821.265 ;
        RECT 1623.040 58.655 1670.640 821.265 ;
        RECT 1673.040 58.655 1720.640 821.265 ;
        RECT 1723.040 58.655 1770.640 821.265 ;
        RECT 1773.040 58.655 1820.640 821.265 ;
        RECT 1823.040 58.655 1870.640 821.265 ;
        RECT 1873.040 58.655 1920.640 821.265 ;
        RECT 1923.040 58.655 1970.640 821.265 ;
        RECT 1973.040 58.655 2014.505 821.265 ;
  END
END pwm_top
END LIBRARY

