magic
tech sky130A
magscale 1 2
timestamp 1647668502
<< obsli1 >>
rect 1104 2159 318872 137649
<< obsm1 >>
rect 1104 1096 318872 138032
<< metal2 >>
rect 1398 139200 1454 140000
rect 4158 139200 4214 140000
rect 7010 139200 7066 140000
rect 9770 139200 9826 140000
rect 12622 139200 12678 140000
rect 15382 139200 15438 140000
rect 18234 139200 18290 140000
rect 20994 139200 21050 140000
rect 23846 139200 23902 140000
rect 26606 139200 26662 140000
rect 29458 139200 29514 140000
rect 32218 139200 32274 140000
rect 35070 139200 35126 140000
rect 37830 139200 37886 140000
rect 40682 139200 40738 140000
rect 43442 139200 43498 140000
rect 46294 139200 46350 140000
rect 49054 139200 49110 140000
rect 51906 139200 51962 140000
rect 54666 139200 54722 140000
rect 57518 139200 57574 140000
rect 60278 139200 60334 140000
rect 63130 139200 63186 140000
rect 65890 139200 65946 140000
rect 68742 139200 68798 140000
rect 71502 139200 71558 140000
rect 74354 139200 74410 140000
rect 77114 139200 77170 140000
rect 79966 139200 80022 140000
rect 82726 139200 82782 140000
rect 85578 139200 85634 140000
rect 88338 139200 88394 140000
rect 91190 139200 91246 140000
rect 93950 139200 94006 140000
rect 96802 139200 96858 140000
rect 99562 139200 99618 140000
rect 102414 139200 102470 140000
rect 105174 139200 105230 140000
rect 108026 139200 108082 140000
rect 110786 139200 110842 140000
rect 113638 139200 113694 140000
rect 116398 139200 116454 140000
rect 119250 139200 119306 140000
rect 122010 139200 122066 140000
rect 124862 139200 124918 140000
rect 127622 139200 127678 140000
rect 130474 139200 130530 140000
rect 133234 139200 133290 140000
rect 136086 139200 136142 140000
rect 138846 139200 138902 140000
rect 141698 139200 141754 140000
rect 144458 139200 144514 140000
rect 147310 139200 147366 140000
rect 150070 139200 150126 140000
rect 152922 139200 152978 140000
rect 155682 139200 155738 140000
rect 158534 139200 158590 140000
rect 161386 139200 161442 140000
rect 164146 139200 164202 140000
rect 166998 139200 167054 140000
rect 169758 139200 169814 140000
rect 172610 139200 172666 140000
rect 175370 139200 175426 140000
rect 178222 139200 178278 140000
rect 180982 139200 181038 140000
rect 183834 139200 183890 140000
rect 186594 139200 186650 140000
rect 189446 139200 189502 140000
rect 192206 139200 192262 140000
rect 195058 139200 195114 140000
rect 197818 139200 197874 140000
rect 200670 139200 200726 140000
rect 203430 139200 203486 140000
rect 206282 139200 206338 140000
rect 209042 139200 209098 140000
rect 211894 139200 211950 140000
rect 214654 139200 214710 140000
rect 217506 139200 217562 140000
rect 220266 139200 220322 140000
rect 223118 139200 223174 140000
rect 225878 139200 225934 140000
rect 228730 139200 228786 140000
rect 231490 139200 231546 140000
rect 234342 139200 234398 140000
rect 237102 139200 237158 140000
rect 239954 139200 240010 140000
rect 242714 139200 242770 140000
rect 245566 139200 245622 140000
rect 248326 139200 248382 140000
rect 251178 139200 251234 140000
rect 253938 139200 253994 140000
rect 256790 139200 256846 140000
rect 259550 139200 259606 140000
rect 262402 139200 262458 140000
rect 265162 139200 265218 140000
rect 268014 139200 268070 140000
rect 270774 139200 270830 140000
rect 273626 139200 273682 140000
rect 276386 139200 276442 140000
rect 279238 139200 279294 140000
rect 281998 139200 282054 140000
rect 284850 139200 284906 140000
rect 287610 139200 287666 140000
rect 290462 139200 290518 140000
rect 293222 139200 293278 140000
rect 296074 139200 296130 140000
rect 298834 139200 298890 140000
rect 301686 139200 301742 140000
rect 304446 139200 304502 140000
rect 307298 139200 307354 140000
rect 310058 139200 310114 140000
rect 312910 139200 312966 140000
rect 315670 139200 315726 140000
rect 318522 139200 318578 140000
rect 1398 0 1454 800
rect 4250 0 4306 800
rect 7194 0 7250 800
rect 10138 0 10194 800
rect 13082 0 13138 800
rect 16026 0 16082 800
rect 18970 0 19026 800
rect 21914 0 21970 800
rect 24858 0 24914 800
rect 27802 0 27858 800
rect 30746 0 30802 800
rect 33598 0 33654 800
rect 36542 0 36598 800
rect 39486 0 39542 800
rect 42430 0 42486 800
rect 45374 0 45430 800
rect 48318 0 48374 800
rect 51262 0 51318 800
rect 54206 0 54262 800
rect 57150 0 57206 800
rect 60094 0 60150 800
rect 63038 0 63094 800
rect 65890 0 65946 800
rect 68834 0 68890 800
rect 71778 0 71834 800
rect 74722 0 74778 800
rect 77666 0 77722 800
rect 80610 0 80666 800
rect 83554 0 83610 800
rect 86498 0 86554 800
rect 89442 0 89498 800
rect 92386 0 92442 800
rect 95330 0 95386 800
rect 98182 0 98238 800
rect 101126 0 101182 800
rect 104070 0 104126 800
rect 107014 0 107070 800
rect 109958 0 110014 800
rect 112902 0 112958 800
rect 115846 0 115902 800
rect 118790 0 118846 800
rect 121734 0 121790 800
rect 124678 0 124734 800
rect 127622 0 127678 800
rect 130474 0 130530 800
rect 133418 0 133474 800
rect 136362 0 136418 800
rect 139306 0 139362 800
rect 142250 0 142306 800
rect 145194 0 145250 800
rect 148138 0 148194 800
rect 151082 0 151138 800
rect 154026 0 154082 800
rect 156970 0 157026 800
rect 159914 0 159970 800
rect 162766 0 162822 800
rect 165710 0 165766 800
rect 168654 0 168710 800
rect 171598 0 171654 800
rect 174542 0 174598 800
rect 177486 0 177542 800
rect 180430 0 180486 800
rect 183374 0 183430 800
rect 186318 0 186374 800
rect 189262 0 189318 800
rect 192206 0 192262 800
rect 195058 0 195114 800
rect 198002 0 198058 800
rect 200946 0 201002 800
rect 203890 0 203946 800
rect 206834 0 206890 800
rect 209778 0 209834 800
rect 212722 0 212778 800
rect 215666 0 215722 800
rect 218610 0 218666 800
rect 221554 0 221610 800
rect 224498 0 224554 800
rect 227350 0 227406 800
rect 230294 0 230350 800
rect 233238 0 233294 800
rect 236182 0 236238 800
rect 239126 0 239182 800
rect 242070 0 242126 800
rect 245014 0 245070 800
rect 247958 0 248014 800
rect 250902 0 250958 800
rect 253846 0 253902 800
rect 256790 0 256846 800
rect 259642 0 259698 800
rect 262586 0 262642 800
rect 265530 0 265586 800
rect 268474 0 268530 800
rect 271418 0 271474 800
rect 274362 0 274418 800
rect 277306 0 277362 800
rect 280250 0 280306 800
rect 283194 0 283250 800
rect 286138 0 286194 800
rect 289082 0 289138 800
rect 291934 0 291990 800
rect 294878 0 294934 800
rect 297822 0 297878 800
rect 300766 0 300822 800
rect 303710 0 303766 800
rect 306654 0 306710 800
rect 309598 0 309654 800
rect 312542 0 312598 800
rect 315486 0 315542 800
rect 318430 0 318486 800
<< obsm2 >>
rect 1510 139144 4102 139369
rect 4270 139144 6954 139369
rect 7122 139144 9714 139369
rect 9882 139144 12566 139369
rect 12734 139144 15326 139369
rect 15494 139144 18178 139369
rect 18346 139144 20938 139369
rect 21106 139144 23790 139369
rect 23958 139144 26550 139369
rect 26718 139144 29402 139369
rect 29570 139144 32162 139369
rect 32330 139144 35014 139369
rect 35182 139144 37774 139369
rect 37942 139144 40626 139369
rect 40794 139144 43386 139369
rect 43554 139144 46238 139369
rect 46406 139144 48998 139369
rect 49166 139144 51850 139369
rect 52018 139144 54610 139369
rect 54778 139144 57462 139369
rect 57630 139144 60222 139369
rect 60390 139144 63074 139369
rect 63242 139144 65834 139369
rect 66002 139144 68686 139369
rect 68854 139144 71446 139369
rect 71614 139144 74298 139369
rect 74466 139144 77058 139369
rect 77226 139144 79910 139369
rect 80078 139144 82670 139369
rect 82838 139144 85522 139369
rect 85690 139144 88282 139369
rect 88450 139144 91134 139369
rect 91302 139144 93894 139369
rect 94062 139144 96746 139369
rect 96914 139144 99506 139369
rect 99674 139144 102358 139369
rect 102526 139144 105118 139369
rect 105286 139144 107970 139369
rect 108138 139144 110730 139369
rect 110898 139144 113582 139369
rect 113750 139144 116342 139369
rect 116510 139144 119194 139369
rect 119362 139144 121954 139369
rect 122122 139144 124806 139369
rect 124974 139144 127566 139369
rect 127734 139144 130418 139369
rect 130586 139144 133178 139369
rect 133346 139144 136030 139369
rect 136198 139144 138790 139369
rect 138958 139144 141642 139369
rect 141810 139144 144402 139369
rect 144570 139144 147254 139369
rect 147422 139144 150014 139369
rect 150182 139144 152866 139369
rect 153034 139144 155626 139369
rect 155794 139144 158478 139369
rect 158646 139144 161330 139369
rect 161498 139144 164090 139369
rect 164258 139144 166942 139369
rect 167110 139144 169702 139369
rect 169870 139144 172554 139369
rect 172722 139144 175314 139369
rect 175482 139144 178166 139369
rect 178334 139144 180926 139369
rect 181094 139144 183778 139369
rect 183946 139144 186538 139369
rect 186706 139144 189390 139369
rect 189558 139144 192150 139369
rect 192318 139144 195002 139369
rect 195170 139144 197762 139369
rect 197930 139144 200614 139369
rect 200782 139144 203374 139369
rect 203542 139144 206226 139369
rect 206394 139144 208986 139369
rect 209154 139144 211838 139369
rect 212006 139144 214598 139369
rect 214766 139144 217450 139369
rect 217618 139144 220210 139369
rect 220378 139144 223062 139369
rect 223230 139144 225822 139369
rect 225990 139144 228674 139369
rect 228842 139144 231434 139369
rect 231602 139144 234286 139369
rect 234454 139144 237046 139369
rect 237214 139144 239898 139369
rect 240066 139144 242658 139369
rect 242826 139144 245510 139369
rect 245678 139144 248270 139369
rect 248438 139144 251122 139369
rect 251290 139144 253882 139369
rect 254050 139144 256734 139369
rect 256902 139144 259494 139369
rect 259662 139144 262346 139369
rect 262514 139144 265106 139369
rect 265274 139144 267958 139369
rect 268126 139144 270718 139369
rect 270886 139144 273570 139369
rect 273738 139144 276330 139369
rect 276498 139144 279182 139369
rect 279350 139144 281942 139369
rect 282110 139144 284794 139369
rect 284962 139144 287554 139369
rect 287722 139144 290406 139369
rect 290574 139144 293166 139369
rect 293334 139144 296018 139369
rect 296186 139144 298778 139369
rect 298946 139144 301630 139369
rect 301798 139144 304390 139369
rect 304558 139144 307242 139369
rect 307410 139144 310002 139369
rect 310170 139144 312854 139369
rect 313022 139144 315614 139369
rect 315782 139144 318466 139369
rect 1400 856 318522 139144
rect 1510 575 4194 856
rect 4362 575 7138 856
rect 7306 575 10082 856
rect 10250 575 13026 856
rect 13194 575 15970 856
rect 16138 575 18914 856
rect 19082 575 21858 856
rect 22026 575 24802 856
rect 24970 575 27746 856
rect 27914 575 30690 856
rect 30858 575 33542 856
rect 33710 575 36486 856
rect 36654 575 39430 856
rect 39598 575 42374 856
rect 42542 575 45318 856
rect 45486 575 48262 856
rect 48430 575 51206 856
rect 51374 575 54150 856
rect 54318 575 57094 856
rect 57262 575 60038 856
rect 60206 575 62982 856
rect 63150 575 65834 856
rect 66002 575 68778 856
rect 68946 575 71722 856
rect 71890 575 74666 856
rect 74834 575 77610 856
rect 77778 575 80554 856
rect 80722 575 83498 856
rect 83666 575 86442 856
rect 86610 575 89386 856
rect 89554 575 92330 856
rect 92498 575 95274 856
rect 95442 575 98126 856
rect 98294 575 101070 856
rect 101238 575 104014 856
rect 104182 575 106958 856
rect 107126 575 109902 856
rect 110070 575 112846 856
rect 113014 575 115790 856
rect 115958 575 118734 856
rect 118902 575 121678 856
rect 121846 575 124622 856
rect 124790 575 127566 856
rect 127734 575 130418 856
rect 130586 575 133362 856
rect 133530 575 136306 856
rect 136474 575 139250 856
rect 139418 575 142194 856
rect 142362 575 145138 856
rect 145306 575 148082 856
rect 148250 575 151026 856
rect 151194 575 153970 856
rect 154138 575 156914 856
rect 157082 575 159858 856
rect 160026 575 162710 856
rect 162878 575 165654 856
rect 165822 575 168598 856
rect 168766 575 171542 856
rect 171710 575 174486 856
rect 174654 575 177430 856
rect 177598 575 180374 856
rect 180542 575 183318 856
rect 183486 575 186262 856
rect 186430 575 189206 856
rect 189374 575 192150 856
rect 192318 575 195002 856
rect 195170 575 197946 856
rect 198114 575 200890 856
rect 201058 575 203834 856
rect 204002 575 206778 856
rect 206946 575 209722 856
rect 209890 575 212666 856
rect 212834 575 215610 856
rect 215778 575 218554 856
rect 218722 575 221498 856
rect 221666 575 224442 856
rect 224610 575 227294 856
rect 227462 575 230238 856
rect 230406 575 233182 856
rect 233350 575 236126 856
rect 236294 575 239070 856
rect 239238 575 242014 856
rect 242182 575 244958 856
rect 245126 575 247902 856
rect 248070 575 250846 856
rect 251014 575 253790 856
rect 253958 575 256734 856
rect 256902 575 259586 856
rect 259754 575 262530 856
rect 262698 575 265474 856
rect 265642 575 268418 856
rect 268586 575 271362 856
rect 271530 575 274306 856
rect 274474 575 277250 856
rect 277418 575 280194 856
rect 280362 575 283138 856
rect 283306 575 286082 856
rect 286250 575 289026 856
rect 289194 575 291878 856
rect 292046 575 294822 856
rect 294990 575 297766 856
rect 297934 575 300710 856
rect 300878 575 303654 856
rect 303822 575 306598 856
rect 306766 575 309542 856
rect 309710 575 312486 856
rect 312654 575 315430 856
rect 315598 575 318374 856
<< metal3 >>
rect 0 139544 800 139664
rect 319200 139272 320000 139392
rect 0 139000 800 139120
rect 0 138456 800 138576
rect 319200 138184 320000 138304
rect 0 137912 800 138032
rect 0 137368 800 137488
rect 319200 137096 320000 137216
rect 0 136824 800 136944
rect 0 136280 800 136400
rect 319200 136008 320000 136128
rect 0 135736 800 135856
rect 0 135192 800 135312
rect 319200 134920 320000 135040
rect 0 134648 800 134768
rect 0 134104 800 134224
rect 319200 133832 320000 133952
rect 0 133560 800 133680
rect 0 133016 800 133136
rect 319200 132744 320000 132864
rect 0 132472 800 132592
rect 0 131928 800 132048
rect 319200 131656 320000 131776
rect 0 131384 800 131504
rect 0 130840 800 130960
rect 319200 130568 320000 130688
rect 0 130296 800 130416
rect 0 129752 800 129872
rect 319200 129480 320000 129600
rect 0 129208 800 129328
rect 0 128664 800 128784
rect 319200 128392 320000 128512
rect 0 128120 800 128240
rect 0 127576 800 127696
rect 319200 127304 320000 127424
rect 0 127032 800 127152
rect 0 126488 800 126608
rect 319200 126216 320000 126336
rect 0 125944 800 126064
rect 0 125400 800 125520
rect 319200 125128 320000 125248
rect 0 124856 800 124976
rect 0 124312 800 124432
rect 319200 124040 320000 124160
rect 0 123768 800 123888
rect 0 123224 800 123344
rect 319200 122952 320000 123072
rect 0 122680 800 122800
rect 0 122136 800 122256
rect 319200 121864 320000 121984
rect 0 121592 800 121712
rect 0 121048 800 121168
rect 319200 120776 320000 120896
rect 0 120504 800 120624
rect 0 119960 800 120080
rect 319200 119688 320000 119808
rect 0 119416 800 119536
rect 0 118872 800 118992
rect 319200 118600 320000 118720
rect 0 118328 800 118448
rect 0 117784 800 117904
rect 319200 117512 320000 117632
rect 0 117240 800 117360
rect 0 116696 800 116816
rect 319200 116424 320000 116544
rect 0 116152 800 116272
rect 0 115608 800 115728
rect 319200 115336 320000 115456
rect 0 115064 800 115184
rect 0 114520 800 114640
rect 319200 114248 320000 114368
rect 0 113976 800 114096
rect 0 113432 800 113552
rect 319200 113160 320000 113280
rect 0 112888 800 113008
rect 0 112344 800 112464
rect 319200 111936 320000 112056
rect 0 111664 800 111784
rect 0 111120 800 111240
rect 319200 110848 320000 110968
rect 0 110576 800 110696
rect 0 110032 800 110152
rect 319200 109760 320000 109880
rect 0 109488 800 109608
rect 0 108944 800 109064
rect 319200 108672 320000 108792
rect 0 108400 800 108520
rect 0 107856 800 107976
rect 319200 107584 320000 107704
rect 0 107312 800 107432
rect 0 106768 800 106888
rect 319200 106496 320000 106616
rect 0 106224 800 106344
rect 0 105680 800 105800
rect 319200 105408 320000 105528
rect 0 105136 800 105256
rect 0 104592 800 104712
rect 319200 104320 320000 104440
rect 0 104048 800 104168
rect 0 103504 800 103624
rect 319200 103232 320000 103352
rect 0 102960 800 103080
rect 0 102416 800 102536
rect 319200 102144 320000 102264
rect 0 101872 800 101992
rect 0 101328 800 101448
rect 319200 101056 320000 101176
rect 0 100784 800 100904
rect 0 100240 800 100360
rect 319200 99968 320000 100088
rect 0 99696 800 99816
rect 0 99152 800 99272
rect 319200 98880 320000 99000
rect 0 98608 800 98728
rect 0 98064 800 98184
rect 319200 97792 320000 97912
rect 0 97520 800 97640
rect 0 96976 800 97096
rect 319200 96704 320000 96824
rect 0 96432 800 96552
rect 0 95888 800 96008
rect 319200 95616 320000 95736
rect 0 95344 800 95464
rect 0 94800 800 94920
rect 319200 94528 320000 94648
rect 0 94256 800 94376
rect 0 93712 800 93832
rect 319200 93440 320000 93560
rect 0 93168 800 93288
rect 0 92624 800 92744
rect 319200 92352 320000 92472
rect 0 92080 800 92200
rect 0 91536 800 91656
rect 319200 91264 320000 91384
rect 0 90992 800 91112
rect 0 90448 800 90568
rect 319200 90176 320000 90296
rect 0 89904 800 90024
rect 0 89360 800 89480
rect 319200 89088 320000 89208
rect 0 88816 800 88936
rect 0 88272 800 88392
rect 319200 88000 320000 88120
rect 0 87728 800 87848
rect 0 87184 800 87304
rect 319200 86912 320000 87032
rect 0 86640 800 86760
rect 0 86096 800 86216
rect 319200 85824 320000 85944
rect 0 85552 800 85672
rect 0 85008 800 85128
rect 319200 84736 320000 84856
rect 0 84464 800 84584
rect 0 83784 800 83904
rect 319200 83512 320000 83632
rect 0 83240 800 83360
rect 0 82696 800 82816
rect 319200 82424 320000 82544
rect 0 82152 800 82272
rect 0 81608 800 81728
rect 319200 81336 320000 81456
rect 0 81064 800 81184
rect 0 80520 800 80640
rect 319200 80248 320000 80368
rect 0 79976 800 80096
rect 0 79432 800 79552
rect 319200 79160 320000 79280
rect 0 78888 800 79008
rect 0 78344 800 78464
rect 319200 78072 320000 78192
rect 0 77800 800 77920
rect 0 77256 800 77376
rect 319200 76984 320000 77104
rect 0 76712 800 76832
rect 0 76168 800 76288
rect 319200 75896 320000 76016
rect 0 75624 800 75744
rect 0 75080 800 75200
rect 319200 74808 320000 74928
rect 0 74536 800 74656
rect 0 73992 800 74112
rect 319200 73720 320000 73840
rect 0 73448 800 73568
rect 0 72904 800 73024
rect 319200 72632 320000 72752
rect 0 72360 800 72480
rect 0 71816 800 71936
rect 319200 71544 320000 71664
rect 0 71272 800 71392
rect 0 70728 800 70848
rect 319200 70456 320000 70576
rect 0 70184 800 70304
rect 0 69640 800 69760
rect 319200 69368 320000 69488
rect 0 69096 800 69216
rect 0 68552 800 68672
rect 319200 68280 320000 68400
rect 0 68008 800 68128
rect 0 67464 800 67584
rect 319200 67192 320000 67312
rect 0 66920 800 67040
rect 0 66376 800 66496
rect 319200 66104 320000 66224
rect 0 65832 800 65952
rect 0 65288 800 65408
rect 319200 65016 320000 65136
rect 0 64744 800 64864
rect 0 64200 800 64320
rect 319200 63928 320000 64048
rect 0 63656 800 63776
rect 0 63112 800 63232
rect 319200 62840 320000 62960
rect 0 62568 800 62688
rect 0 62024 800 62144
rect 319200 61752 320000 61872
rect 0 61480 800 61600
rect 0 60936 800 61056
rect 319200 60664 320000 60784
rect 0 60392 800 60512
rect 0 59848 800 59968
rect 319200 59576 320000 59696
rect 0 59304 800 59424
rect 0 58760 800 58880
rect 319200 58488 320000 58608
rect 0 58216 800 58336
rect 0 57672 800 57792
rect 319200 57400 320000 57520
rect 0 57128 800 57248
rect 0 56584 800 56704
rect 319200 56176 320000 56296
rect 0 55904 800 56024
rect 0 55360 800 55480
rect 319200 55088 320000 55208
rect 0 54816 800 54936
rect 0 54272 800 54392
rect 319200 54000 320000 54120
rect 0 53728 800 53848
rect 0 53184 800 53304
rect 319200 52912 320000 53032
rect 0 52640 800 52760
rect 0 52096 800 52216
rect 319200 51824 320000 51944
rect 0 51552 800 51672
rect 0 51008 800 51128
rect 319200 50736 320000 50856
rect 0 50464 800 50584
rect 0 49920 800 50040
rect 319200 49648 320000 49768
rect 0 49376 800 49496
rect 0 48832 800 48952
rect 319200 48560 320000 48680
rect 0 48288 800 48408
rect 0 47744 800 47864
rect 319200 47472 320000 47592
rect 0 47200 800 47320
rect 0 46656 800 46776
rect 319200 46384 320000 46504
rect 0 46112 800 46232
rect 0 45568 800 45688
rect 319200 45296 320000 45416
rect 0 45024 800 45144
rect 0 44480 800 44600
rect 319200 44208 320000 44328
rect 0 43936 800 44056
rect 0 43392 800 43512
rect 319200 43120 320000 43240
rect 0 42848 800 42968
rect 0 42304 800 42424
rect 319200 42032 320000 42152
rect 0 41760 800 41880
rect 0 41216 800 41336
rect 319200 40944 320000 41064
rect 0 40672 800 40792
rect 0 40128 800 40248
rect 319200 39856 320000 39976
rect 0 39584 800 39704
rect 0 39040 800 39160
rect 319200 38768 320000 38888
rect 0 38496 800 38616
rect 0 37952 800 38072
rect 319200 37680 320000 37800
rect 0 37408 800 37528
rect 0 36864 800 36984
rect 319200 36592 320000 36712
rect 0 36320 800 36440
rect 0 35776 800 35896
rect 319200 35504 320000 35624
rect 0 35232 800 35352
rect 0 34688 800 34808
rect 319200 34416 320000 34536
rect 0 34144 800 34264
rect 0 33600 800 33720
rect 319200 33328 320000 33448
rect 0 33056 800 33176
rect 0 32512 800 32632
rect 319200 32240 320000 32360
rect 0 31968 800 32088
rect 0 31424 800 31544
rect 319200 31152 320000 31272
rect 0 30880 800 31000
rect 0 30336 800 30456
rect 319200 30064 320000 30184
rect 0 29792 800 29912
rect 0 29248 800 29368
rect 319200 28976 320000 29096
rect 0 28704 800 28824
rect 0 28024 800 28144
rect 319200 27752 320000 27872
rect 0 27480 800 27600
rect 0 26936 800 27056
rect 319200 26664 320000 26784
rect 0 26392 800 26512
rect 0 25848 800 25968
rect 319200 25576 320000 25696
rect 0 25304 800 25424
rect 0 24760 800 24880
rect 319200 24488 320000 24608
rect 0 24216 800 24336
rect 0 23672 800 23792
rect 319200 23400 320000 23520
rect 0 23128 800 23248
rect 0 22584 800 22704
rect 319200 22312 320000 22432
rect 0 22040 800 22160
rect 0 21496 800 21616
rect 319200 21224 320000 21344
rect 0 20952 800 21072
rect 0 20408 800 20528
rect 319200 20136 320000 20256
rect 0 19864 800 19984
rect 0 19320 800 19440
rect 319200 19048 320000 19168
rect 0 18776 800 18896
rect 0 18232 800 18352
rect 319200 17960 320000 18080
rect 0 17688 800 17808
rect 0 17144 800 17264
rect 319200 16872 320000 16992
rect 0 16600 800 16720
rect 0 16056 800 16176
rect 319200 15784 320000 15904
rect 0 15512 800 15632
rect 0 14968 800 15088
rect 319200 14696 320000 14816
rect 0 14424 800 14544
rect 0 13880 800 14000
rect 319200 13608 320000 13728
rect 0 13336 800 13456
rect 0 12792 800 12912
rect 319200 12520 320000 12640
rect 0 12248 800 12368
rect 0 11704 800 11824
rect 319200 11432 320000 11552
rect 0 11160 800 11280
rect 0 10616 800 10736
rect 319200 10344 320000 10464
rect 0 10072 800 10192
rect 0 9528 800 9648
rect 319200 9256 320000 9376
rect 0 8984 800 9104
rect 0 8440 800 8560
rect 319200 8168 320000 8288
rect 0 7896 800 8016
rect 0 7352 800 7472
rect 319200 7080 320000 7200
rect 0 6808 800 6928
rect 0 6264 800 6384
rect 319200 5992 320000 6112
rect 0 5720 800 5840
rect 0 5176 800 5296
rect 319200 4904 320000 5024
rect 0 4632 800 4752
rect 0 4088 800 4208
rect 319200 3816 320000 3936
rect 0 3544 800 3664
rect 0 3000 800 3120
rect 319200 2728 320000 2848
rect 0 2456 800 2576
rect 0 1912 800 2032
rect 319200 1640 320000 1760
rect 0 1368 800 1488
rect 0 824 800 944
rect 319200 552 320000 672
rect 0 280 800 400
<< obsm3 >>
rect 2129 139192 319120 139365
rect 2129 138384 319200 139192
rect 2129 138104 319120 138384
rect 2129 137296 319200 138104
rect 2129 137016 319120 137296
rect 2129 136208 319200 137016
rect 2129 135928 319120 136208
rect 2129 135120 319200 135928
rect 2129 134840 319120 135120
rect 2129 134032 319200 134840
rect 2129 133752 319120 134032
rect 2129 132944 319200 133752
rect 2129 132664 319120 132944
rect 2129 131856 319200 132664
rect 2129 131576 319120 131856
rect 2129 130768 319200 131576
rect 2129 130488 319120 130768
rect 2129 129680 319200 130488
rect 2129 129400 319120 129680
rect 2129 128592 319200 129400
rect 2129 128312 319120 128592
rect 2129 127504 319200 128312
rect 2129 127224 319120 127504
rect 2129 126416 319200 127224
rect 2129 126136 319120 126416
rect 2129 125328 319200 126136
rect 2129 125048 319120 125328
rect 2129 124240 319200 125048
rect 2129 123960 319120 124240
rect 2129 123152 319200 123960
rect 2129 122872 319120 123152
rect 2129 122064 319200 122872
rect 2129 121784 319120 122064
rect 2129 120976 319200 121784
rect 2129 120696 319120 120976
rect 2129 119888 319200 120696
rect 2129 119608 319120 119888
rect 2129 118800 319200 119608
rect 2129 118520 319120 118800
rect 2129 117712 319200 118520
rect 2129 117432 319120 117712
rect 2129 116624 319200 117432
rect 2129 116344 319120 116624
rect 2129 115536 319200 116344
rect 2129 115256 319120 115536
rect 2129 114448 319200 115256
rect 2129 114168 319120 114448
rect 2129 113360 319200 114168
rect 2129 113080 319120 113360
rect 2129 112136 319200 113080
rect 2129 111856 319120 112136
rect 2129 111048 319200 111856
rect 2129 110768 319120 111048
rect 2129 109960 319200 110768
rect 2129 109680 319120 109960
rect 2129 108872 319200 109680
rect 2129 108592 319120 108872
rect 2129 107784 319200 108592
rect 2129 107504 319120 107784
rect 2129 106696 319200 107504
rect 2129 106416 319120 106696
rect 2129 105608 319200 106416
rect 2129 105328 319120 105608
rect 2129 104520 319200 105328
rect 2129 104240 319120 104520
rect 2129 103432 319200 104240
rect 2129 103152 319120 103432
rect 2129 102344 319200 103152
rect 2129 102064 319120 102344
rect 2129 101256 319200 102064
rect 2129 100976 319120 101256
rect 2129 100168 319200 100976
rect 2129 99888 319120 100168
rect 2129 99080 319200 99888
rect 2129 98800 319120 99080
rect 2129 97992 319200 98800
rect 2129 97712 319120 97992
rect 2129 96904 319200 97712
rect 2129 96624 319120 96904
rect 2129 95816 319200 96624
rect 2129 95536 319120 95816
rect 2129 94728 319200 95536
rect 2129 94448 319120 94728
rect 2129 93640 319200 94448
rect 2129 93360 319120 93640
rect 2129 92552 319200 93360
rect 2129 92272 319120 92552
rect 2129 91464 319200 92272
rect 2129 91184 319120 91464
rect 2129 90376 319200 91184
rect 2129 90096 319120 90376
rect 2129 89288 319200 90096
rect 2129 89008 319120 89288
rect 2129 88200 319200 89008
rect 2129 87920 319120 88200
rect 2129 87112 319200 87920
rect 2129 86832 319120 87112
rect 2129 86024 319200 86832
rect 2129 85744 319120 86024
rect 2129 84936 319200 85744
rect 2129 84656 319120 84936
rect 2129 83712 319200 84656
rect 2129 83432 319120 83712
rect 2129 82624 319200 83432
rect 2129 82344 319120 82624
rect 2129 81536 319200 82344
rect 2129 81256 319120 81536
rect 2129 80448 319200 81256
rect 2129 80168 319120 80448
rect 2129 79360 319200 80168
rect 2129 79080 319120 79360
rect 2129 78272 319200 79080
rect 2129 77992 319120 78272
rect 2129 77184 319200 77992
rect 2129 76904 319120 77184
rect 2129 76096 319200 76904
rect 2129 75816 319120 76096
rect 2129 75008 319200 75816
rect 2129 74728 319120 75008
rect 2129 73920 319200 74728
rect 2129 73640 319120 73920
rect 2129 72832 319200 73640
rect 2129 72552 319120 72832
rect 2129 71744 319200 72552
rect 2129 71464 319120 71744
rect 2129 70656 319200 71464
rect 2129 70376 319120 70656
rect 2129 69568 319200 70376
rect 2129 69288 319120 69568
rect 2129 68480 319200 69288
rect 2129 68200 319120 68480
rect 2129 67392 319200 68200
rect 2129 67112 319120 67392
rect 2129 66304 319200 67112
rect 2129 66024 319120 66304
rect 2129 65216 319200 66024
rect 2129 64936 319120 65216
rect 2129 64128 319200 64936
rect 2129 63848 319120 64128
rect 2129 63040 319200 63848
rect 2129 62760 319120 63040
rect 2129 61952 319200 62760
rect 2129 61672 319120 61952
rect 2129 60864 319200 61672
rect 2129 60584 319120 60864
rect 2129 59776 319200 60584
rect 2129 59496 319120 59776
rect 2129 58688 319200 59496
rect 2129 58408 319120 58688
rect 2129 57600 319200 58408
rect 2129 57320 319120 57600
rect 2129 56376 319200 57320
rect 2129 56096 319120 56376
rect 2129 55288 319200 56096
rect 2129 55008 319120 55288
rect 2129 54200 319200 55008
rect 2129 53920 319120 54200
rect 2129 53112 319200 53920
rect 2129 52832 319120 53112
rect 2129 52024 319200 52832
rect 2129 51744 319120 52024
rect 2129 50936 319200 51744
rect 2129 50656 319120 50936
rect 2129 49848 319200 50656
rect 2129 49568 319120 49848
rect 2129 48760 319200 49568
rect 2129 48480 319120 48760
rect 2129 47672 319200 48480
rect 2129 47392 319120 47672
rect 2129 46584 319200 47392
rect 2129 46304 319120 46584
rect 2129 45496 319200 46304
rect 2129 45216 319120 45496
rect 2129 44408 319200 45216
rect 2129 44128 319120 44408
rect 2129 43320 319200 44128
rect 2129 43040 319120 43320
rect 2129 42232 319200 43040
rect 2129 41952 319120 42232
rect 2129 41144 319200 41952
rect 2129 40864 319120 41144
rect 2129 40056 319200 40864
rect 2129 39776 319120 40056
rect 2129 38968 319200 39776
rect 2129 38688 319120 38968
rect 2129 37880 319200 38688
rect 2129 37600 319120 37880
rect 2129 36792 319200 37600
rect 2129 36512 319120 36792
rect 2129 35704 319200 36512
rect 2129 35424 319120 35704
rect 2129 34616 319200 35424
rect 2129 34336 319120 34616
rect 2129 33528 319200 34336
rect 2129 33248 319120 33528
rect 2129 32440 319200 33248
rect 2129 32160 319120 32440
rect 2129 31352 319200 32160
rect 2129 31072 319120 31352
rect 2129 30264 319200 31072
rect 2129 29984 319120 30264
rect 2129 29176 319200 29984
rect 2129 28896 319120 29176
rect 2129 27952 319200 28896
rect 2129 27672 319120 27952
rect 2129 26864 319200 27672
rect 2129 26584 319120 26864
rect 2129 25776 319200 26584
rect 2129 25496 319120 25776
rect 2129 24688 319200 25496
rect 2129 24408 319120 24688
rect 2129 23600 319200 24408
rect 2129 23320 319120 23600
rect 2129 22512 319200 23320
rect 2129 22232 319120 22512
rect 2129 21424 319200 22232
rect 2129 21144 319120 21424
rect 2129 20336 319200 21144
rect 2129 20056 319120 20336
rect 2129 19248 319200 20056
rect 2129 18968 319120 19248
rect 2129 18160 319200 18968
rect 2129 17880 319120 18160
rect 2129 17072 319200 17880
rect 2129 16792 319120 17072
rect 2129 15984 319200 16792
rect 2129 15704 319120 15984
rect 2129 14896 319200 15704
rect 2129 14616 319120 14896
rect 2129 13808 319200 14616
rect 2129 13528 319120 13808
rect 2129 12720 319200 13528
rect 2129 12440 319120 12720
rect 2129 11632 319200 12440
rect 2129 11352 319120 11632
rect 2129 10544 319200 11352
rect 2129 10264 319120 10544
rect 2129 9456 319200 10264
rect 2129 9176 319120 9456
rect 2129 8368 319200 9176
rect 2129 8088 319120 8368
rect 2129 7280 319200 8088
rect 2129 7000 319120 7280
rect 2129 6192 319200 7000
rect 2129 5912 319120 6192
rect 2129 5104 319200 5912
rect 2129 4824 319120 5104
rect 2129 4016 319200 4824
rect 2129 3736 319120 4016
rect 2129 2928 319200 3736
rect 2129 2648 319120 2928
rect 2129 1840 319200 2648
rect 2129 1560 319120 1840
rect 2129 752 319200 1560
rect 2129 579 319120 752
<< metal4 >>
rect 4208 2128 4528 137680
rect 14208 2128 14528 137680
rect 24208 2128 24528 137680
rect 34208 2128 34528 137680
rect 44208 2128 44528 137680
rect 54208 2128 54528 137680
rect 64208 2128 64528 137680
rect 74208 2128 74528 137680
rect 84208 2128 84528 137680
rect 94208 2128 94528 137680
rect 104208 2128 104528 137680
rect 114208 2128 114528 137680
rect 124208 2128 124528 137680
rect 134208 2128 134528 137680
rect 144208 2128 144528 137680
rect 154208 2128 154528 137680
rect 164208 2128 164528 137680
rect 174208 2128 174528 137680
rect 184208 2128 184528 137680
rect 194208 2128 194528 137680
rect 204208 2128 204528 137680
rect 214208 2128 214528 137680
rect 224208 2128 224528 137680
rect 234208 2128 234528 137680
rect 244208 2128 244528 137680
rect 254208 2128 254528 137680
rect 264208 2128 264528 137680
rect 274208 2128 274528 137680
rect 284208 2128 284528 137680
rect 294208 2128 294528 137680
rect 304208 2128 304528 137680
rect 314208 2128 314528 137680
<< obsm4 >>
rect 37779 137760 290109 138277
rect 37779 2347 44128 137760
rect 44608 2347 54128 137760
rect 54608 2347 64128 137760
rect 64608 2347 74128 137760
rect 74608 2347 84128 137760
rect 84608 2347 94128 137760
rect 94608 2347 104128 137760
rect 104608 2347 114128 137760
rect 114608 2347 124128 137760
rect 124608 2347 134128 137760
rect 134608 2347 144128 137760
rect 144608 2347 154128 137760
rect 154608 2347 164128 137760
rect 164608 2347 174128 137760
rect 174608 2347 184128 137760
rect 184608 2347 194128 137760
rect 194608 2347 204128 137760
rect 204608 2347 214128 137760
rect 214608 2347 224128 137760
rect 224608 2347 234128 137760
rect 234608 2347 244128 137760
rect 244608 2347 254128 137760
rect 254608 2347 264128 137760
rect 264608 2347 274128 137760
rect 274608 2347 284128 137760
rect 284608 2347 290109 137760
<< labels >>
rlabel metal2 s 1398 139200 1454 140000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 85578 139200 85634 140000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 93950 139200 94006 140000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 102414 139200 102470 140000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 110786 139200 110842 140000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 119250 139200 119306 140000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 127622 139200 127678 140000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 136086 139200 136142 140000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 144458 139200 144514 140000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 152922 139200 152978 140000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 161386 139200 161442 140000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 9770 139200 9826 140000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 169758 139200 169814 140000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 178222 139200 178278 140000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 186594 139200 186650 140000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 195058 139200 195114 140000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 203430 139200 203486 140000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 211894 139200 211950 140000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 220266 139200 220322 140000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 228730 139200 228786 140000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 237102 139200 237158 140000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 245566 139200 245622 140000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 18234 139200 18290 140000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 253938 139200 253994 140000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 262402 139200 262458 140000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 270774 139200 270830 140000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 279238 139200 279294 140000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 287610 139200 287666 140000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 296074 139200 296130 140000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 304446 139200 304502 140000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 312910 139200 312966 140000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 26606 139200 26662 140000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 35070 139200 35126 140000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 43442 139200 43498 140000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 51906 139200 51962 140000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 60278 139200 60334 140000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 68742 139200 68798 140000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 77114 139200 77170 140000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 4158 139200 4214 140000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 88338 139200 88394 140000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 96802 139200 96858 140000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 105174 139200 105230 140000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 113638 139200 113694 140000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 122010 139200 122066 140000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 130474 139200 130530 140000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 138846 139200 138902 140000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 147310 139200 147366 140000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 155682 139200 155738 140000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 164146 139200 164202 140000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 12622 139200 12678 140000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 172610 139200 172666 140000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 180982 139200 181038 140000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 189446 139200 189502 140000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 197818 139200 197874 140000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 206282 139200 206338 140000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 214654 139200 214710 140000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 223118 139200 223174 140000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 231490 139200 231546 140000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 239954 139200 240010 140000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 248326 139200 248382 140000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 20994 139200 21050 140000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 256790 139200 256846 140000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 265162 139200 265218 140000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 273626 139200 273682 140000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 281998 139200 282054 140000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 290462 139200 290518 140000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 298834 139200 298890 140000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 307298 139200 307354 140000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 315670 139200 315726 140000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 29458 139200 29514 140000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 37830 139200 37886 140000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 46294 139200 46350 140000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 54666 139200 54722 140000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 63130 139200 63186 140000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 71502 139200 71558 140000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 79966 139200 80022 140000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 7010 139200 7066 140000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 91190 139200 91246 140000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 99562 139200 99618 140000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 108026 139200 108082 140000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 116398 139200 116454 140000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 124862 139200 124918 140000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 133234 139200 133290 140000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 141698 139200 141754 140000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 150070 139200 150126 140000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 158534 139200 158590 140000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 166998 139200 167054 140000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 15382 139200 15438 140000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 175370 139200 175426 140000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 183834 139200 183890 140000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 192206 139200 192262 140000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 200670 139200 200726 140000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 209042 139200 209098 140000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 217506 139200 217562 140000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 225878 139200 225934 140000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 234342 139200 234398 140000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 242714 139200 242770 140000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 251178 139200 251234 140000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 23846 139200 23902 140000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 259550 139200 259606 140000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 268014 139200 268070 140000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 276386 139200 276442 140000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 284850 139200 284906 140000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 293222 139200 293278 140000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 301686 139200 301742 140000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 310058 139200 310114 140000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 318522 139200 318578 140000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 32218 139200 32274 140000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 40682 139200 40738 140000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 49054 139200 49110 140000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 57518 139200 57574 140000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 65890 139200 65946 140000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 74354 139200 74410 140000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 82726 139200 82782 140000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 312542 0 312598 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 315486 0 315542 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 318430 0 318486 800 6 irq[2]
port 117 nsew signal output
rlabel metal3 s 0 280 800 400 6 la_data_in[0]
port 118 nsew signal input
rlabel metal3 s 0 54816 800 54936 6 la_data_in[100]
port 119 nsew signal input
rlabel metal3 s 0 55360 800 55480 6 la_data_in[101]
port 120 nsew signal input
rlabel metal3 s 0 55904 800 56024 6 la_data_in[102]
port 121 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 la_data_in[103]
port 122 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 la_data_in[104]
port 123 nsew signal input
rlabel metal3 s 0 57672 800 57792 6 la_data_in[105]
port 124 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 la_data_in[106]
port 125 nsew signal input
rlabel metal3 s 0 58760 800 58880 6 la_data_in[107]
port 126 nsew signal input
rlabel metal3 s 0 59304 800 59424 6 la_data_in[108]
port 127 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 la_data_in[109]
port 128 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 la_data_in[10]
port 129 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 la_data_in[110]
port 130 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 la_data_in[111]
port 131 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 la_data_in[112]
port 132 nsew signal input
rlabel metal3 s 0 62024 800 62144 6 la_data_in[113]
port 133 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 la_data_in[114]
port 134 nsew signal input
rlabel metal3 s 0 63112 800 63232 6 la_data_in[115]
port 135 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 la_data_in[116]
port 136 nsew signal input
rlabel metal3 s 0 64200 800 64320 6 la_data_in[117]
port 137 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 la_data_in[118]
port 138 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 la_data_in[119]
port 139 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 la_data_in[11]
port 140 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 la_data_in[120]
port 141 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 la_data_in[121]
port 142 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 la_data_in[122]
port 143 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 la_data_in[123]
port 144 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 la_data_in[124]
port 145 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 la_data_in[125]
port 146 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 la_data_in[126]
port 147 nsew signal input
rlabel metal3 s 0 69640 800 69760 6 la_data_in[127]
port 148 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 la_data_in[12]
port 149 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 la_data_in[13]
port 150 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 la_data_in[14]
port 151 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 la_data_in[15]
port 152 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 la_data_in[16]
port 153 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 la_data_in[17]
port 154 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 la_data_in[18]
port 155 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 la_data_in[19]
port 156 nsew signal input
rlabel metal3 s 0 824 800 944 6 la_data_in[1]
port 157 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 la_data_in[20]
port 158 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 la_data_in[21]
port 159 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 la_data_in[22]
port 160 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 la_data_in[23]
port 161 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 la_data_in[24]
port 162 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 la_data_in[25]
port 163 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 la_data_in[26]
port 164 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 la_data_in[27]
port 165 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 la_data_in[28]
port 166 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 la_data_in[29]
port 167 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 la_data_in[2]
port 168 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 la_data_in[30]
port 169 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 la_data_in[31]
port 170 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 la_data_in[32]
port 171 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 la_data_in[33]
port 172 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 la_data_in[34]
port 173 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 la_data_in[35]
port 174 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 la_data_in[36]
port 175 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 la_data_in[37]
port 176 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 la_data_in[38]
port 177 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 la_data_in[39]
port 178 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 la_data_in[3]
port 179 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 la_data_in[40]
port 180 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 la_data_in[41]
port 181 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 la_data_in[42]
port 182 nsew signal input
rlabel metal3 s 0 23672 800 23792 6 la_data_in[43]
port 183 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 la_data_in[44]
port 184 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 la_data_in[45]
port 185 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 la_data_in[46]
port 186 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 la_data_in[47]
port 187 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 la_data_in[48]
port 188 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 la_data_in[49]
port 189 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 la_data_in[4]
port 190 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 la_data_in[50]
port 191 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 la_data_in[51]
port 192 nsew signal input
rlabel metal3 s 0 28704 800 28824 6 la_data_in[52]
port 193 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 la_data_in[53]
port 194 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 la_data_in[54]
port 195 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 la_data_in[55]
port 196 nsew signal input
rlabel metal3 s 0 30880 800 31000 6 la_data_in[56]
port 197 nsew signal input
rlabel metal3 s 0 31424 800 31544 6 la_data_in[57]
port 198 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 la_data_in[58]
port 199 nsew signal input
rlabel metal3 s 0 32512 800 32632 6 la_data_in[59]
port 200 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 la_data_in[5]
port 201 nsew signal input
rlabel metal3 s 0 33056 800 33176 6 la_data_in[60]
port 202 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 la_data_in[61]
port 203 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 la_data_in[62]
port 204 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 la_data_in[63]
port 205 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 la_data_in[64]
port 206 nsew signal input
rlabel metal3 s 0 35776 800 35896 6 la_data_in[65]
port 207 nsew signal input
rlabel metal3 s 0 36320 800 36440 6 la_data_in[66]
port 208 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 la_data_in[67]
port 209 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 la_data_in[68]
port 210 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 la_data_in[69]
port 211 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 la_data_in[6]
port 212 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 la_data_in[70]
port 213 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 la_data_in[71]
port 214 nsew signal input
rlabel metal3 s 0 39584 800 39704 6 la_data_in[72]
port 215 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 la_data_in[73]
port 216 nsew signal input
rlabel metal3 s 0 40672 800 40792 6 la_data_in[74]
port 217 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 la_data_in[75]
port 218 nsew signal input
rlabel metal3 s 0 41760 800 41880 6 la_data_in[76]
port 219 nsew signal input
rlabel metal3 s 0 42304 800 42424 6 la_data_in[77]
port 220 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 la_data_in[78]
port 221 nsew signal input
rlabel metal3 s 0 43392 800 43512 6 la_data_in[79]
port 222 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 la_data_in[7]
port 223 nsew signal input
rlabel metal3 s 0 43936 800 44056 6 la_data_in[80]
port 224 nsew signal input
rlabel metal3 s 0 44480 800 44600 6 la_data_in[81]
port 225 nsew signal input
rlabel metal3 s 0 45024 800 45144 6 la_data_in[82]
port 226 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 la_data_in[83]
port 227 nsew signal input
rlabel metal3 s 0 46112 800 46232 6 la_data_in[84]
port 228 nsew signal input
rlabel metal3 s 0 46656 800 46776 6 la_data_in[85]
port 229 nsew signal input
rlabel metal3 s 0 47200 800 47320 6 la_data_in[86]
port 230 nsew signal input
rlabel metal3 s 0 47744 800 47864 6 la_data_in[87]
port 231 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 la_data_in[88]
port 232 nsew signal input
rlabel metal3 s 0 48832 800 48952 6 la_data_in[89]
port 233 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 la_data_in[8]
port 234 nsew signal input
rlabel metal3 s 0 49376 800 49496 6 la_data_in[90]
port 235 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 la_data_in[91]
port 236 nsew signal input
rlabel metal3 s 0 50464 800 50584 6 la_data_in[92]
port 237 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 la_data_in[93]
port 238 nsew signal input
rlabel metal3 s 0 51552 800 51672 6 la_data_in[94]
port 239 nsew signal input
rlabel metal3 s 0 52096 800 52216 6 la_data_in[95]
port 240 nsew signal input
rlabel metal3 s 0 52640 800 52760 6 la_data_in[96]
port 241 nsew signal input
rlabel metal3 s 0 53184 800 53304 6 la_data_in[97]
port 242 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 la_data_in[98]
port 243 nsew signal input
rlabel metal3 s 0 54272 800 54392 6 la_data_in[99]
port 244 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 la_data_in[9]
port 245 nsew signal input
rlabel metal3 s 319200 552 320000 672 6 la_data_out[0]
port 246 nsew signal output
rlabel metal3 s 319200 109760 320000 109880 6 la_data_out[100]
port 247 nsew signal output
rlabel metal3 s 319200 110848 320000 110968 6 la_data_out[101]
port 248 nsew signal output
rlabel metal3 s 319200 111936 320000 112056 6 la_data_out[102]
port 249 nsew signal output
rlabel metal3 s 319200 113160 320000 113280 6 la_data_out[103]
port 250 nsew signal output
rlabel metal3 s 319200 114248 320000 114368 6 la_data_out[104]
port 251 nsew signal output
rlabel metal3 s 319200 115336 320000 115456 6 la_data_out[105]
port 252 nsew signal output
rlabel metal3 s 319200 116424 320000 116544 6 la_data_out[106]
port 253 nsew signal output
rlabel metal3 s 319200 117512 320000 117632 6 la_data_out[107]
port 254 nsew signal output
rlabel metal3 s 319200 118600 320000 118720 6 la_data_out[108]
port 255 nsew signal output
rlabel metal3 s 319200 119688 320000 119808 6 la_data_out[109]
port 256 nsew signal output
rlabel metal3 s 319200 11432 320000 11552 6 la_data_out[10]
port 257 nsew signal output
rlabel metal3 s 319200 120776 320000 120896 6 la_data_out[110]
port 258 nsew signal output
rlabel metal3 s 319200 121864 320000 121984 6 la_data_out[111]
port 259 nsew signal output
rlabel metal3 s 319200 122952 320000 123072 6 la_data_out[112]
port 260 nsew signal output
rlabel metal3 s 319200 124040 320000 124160 6 la_data_out[113]
port 261 nsew signal output
rlabel metal3 s 319200 125128 320000 125248 6 la_data_out[114]
port 262 nsew signal output
rlabel metal3 s 319200 126216 320000 126336 6 la_data_out[115]
port 263 nsew signal output
rlabel metal3 s 319200 127304 320000 127424 6 la_data_out[116]
port 264 nsew signal output
rlabel metal3 s 319200 128392 320000 128512 6 la_data_out[117]
port 265 nsew signal output
rlabel metal3 s 319200 129480 320000 129600 6 la_data_out[118]
port 266 nsew signal output
rlabel metal3 s 319200 130568 320000 130688 6 la_data_out[119]
port 267 nsew signal output
rlabel metal3 s 319200 12520 320000 12640 6 la_data_out[11]
port 268 nsew signal output
rlabel metal3 s 319200 131656 320000 131776 6 la_data_out[120]
port 269 nsew signal output
rlabel metal3 s 319200 132744 320000 132864 6 la_data_out[121]
port 270 nsew signal output
rlabel metal3 s 319200 133832 320000 133952 6 la_data_out[122]
port 271 nsew signal output
rlabel metal3 s 319200 134920 320000 135040 6 la_data_out[123]
port 272 nsew signal output
rlabel metal3 s 319200 136008 320000 136128 6 la_data_out[124]
port 273 nsew signal output
rlabel metal3 s 319200 137096 320000 137216 6 la_data_out[125]
port 274 nsew signal output
rlabel metal3 s 319200 138184 320000 138304 6 la_data_out[126]
port 275 nsew signal output
rlabel metal3 s 319200 139272 320000 139392 6 la_data_out[127]
port 276 nsew signal output
rlabel metal3 s 319200 13608 320000 13728 6 la_data_out[12]
port 277 nsew signal output
rlabel metal3 s 319200 14696 320000 14816 6 la_data_out[13]
port 278 nsew signal output
rlabel metal3 s 319200 15784 320000 15904 6 la_data_out[14]
port 279 nsew signal output
rlabel metal3 s 319200 16872 320000 16992 6 la_data_out[15]
port 280 nsew signal output
rlabel metal3 s 319200 17960 320000 18080 6 la_data_out[16]
port 281 nsew signal output
rlabel metal3 s 319200 19048 320000 19168 6 la_data_out[17]
port 282 nsew signal output
rlabel metal3 s 319200 20136 320000 20256 6 la_data_out[18]
port 283 nsew signal output
rlabel metal3 s 319200 21224 320000 21344 6 la_data_out[19]
port 284 nsew signal output
rlabel metal3 s 319200 1640 320000 1760 6 la_data_out[1]
port 285 nsew signal output
rlabel metal3 s 319200 22312 320000 22432 6 la_data_out[20]
port 286 nsew signal output
rlabel metal3 s 319200 23400 320000 23520 6 la_data_out[21]
port 287 nsew signal output
rlabel metal3 s 319200 24488 320000 24608 6 la_data_out[22]
port 288 nsew signal output
rlabel metal3 s 319200 25576 320000 25696 6 la_data_out[23]
port 289 nsew signal output
rlabel metal3 s 319200 26664 320000 26784 6 la_data_out[24]
port 290 nsew signal output
rlabel metal3 s 319200 27752 320000 27872 6 la_data_out[25]
port 291 nsew signal output
rlabel metal3 s 319200 28976 320000 29096 6 la_data_out[26]
port 292 nsew signal output
rlabel metal3 s 319200 30064 320000 30184 6 la_data_out[27]
port 293 nsew signal output
rlabel metal3 s 319200 31152 320000 31272 6 la_data_out[28]
port 294 nsew signal output
rlabel metal3 s 319200 32240 320000 32360 6 la_data_out[29]
port 295 nsew signal output
rlabel metal3 s 319200 2728 320000 2848 6 la_data_out[2]
port 296 nsew signal output
rlabel metal3 s 319200 33328 320000 33448 6 la_data_out[30]
port 297 nsew signal output
rlabel metal3 s 319200 34416 320000 34536 6 la_data_out[31]
port 298 nsew signal output
rlabel metal3 s 319200 35504 320000 35624 6 la_data_out[32]
port 299 nsew signal output
rlabel metal3 s 319200 36592 320000 36712 6 la_data_out[33]
port 300 nsew signal output
rlabel metal3 s 319200 37680 320000 37800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal3 s 319200 38768 320000 38888 6 la_data_out[35]
port 302 nsew signal output
rlabel metal3 s 319200 39856 320000 39976 6 la_data_out[36]
port 303 nsew signal output
rlabel metal3 s 319200 40944 320000 41064 6 la_data_out[37]
port 304 nsew signal output
rlabel metal3 s 319200 42032 320000 42152 6 la_data_out[38]
port 305 nsew signal output
rlabel metal3 s 319200 43120 320000 43240 6 la_data_out[39]
port 306 nsew signal output
rlabel metal3 s 319200 3816 320000 3936 6 la_data_out[3]
port 307 nsew signal output
rlabel metal3 s 319200 44208 320000 44328 6 la_data_out[40]
port 308 nsew signal output
rlabel metal3 s 319200 45296 320000 45416 6 la_data_out[41]
port 309 nsew signal output
rlabel metal3 s 319200 46384 320000 46504 6 la_data_out[42]
port 310 nsew signal output
rlabel metal3 s 319200 47472 320000 47592 6 la_data_out[43]
port 311 nsew signal output
rlabel metal3 s 319200 48560 320000 48680 6 la_data_out[44]
port 312 nsew signal output
rlabel metal3 s 319200 49648 320000 49768 6 la_data_out[45]
port 313 nsew signal output
rlabel metal3 s 319200 50736 320000 50856 6 la_data_out[46]
port 314 nsew signal output
rlabel metal3 s 319200 51824 320000 51944 6 la_data_out[47]
port 315 nsew signal output
rlabel metal3 s 319200 52912 320000 53032 6 la_data_out[48]
port 316 nsew signal output
rlabel metal3 s 319200 54000 320000 54120 6 la_data_out[49]
port 317 nsew signal output
rlabel metal3 s 319200 4904 320000 5024 6 la_data_out[4]
port 318 nsew signal output
rlabel metal3 s 319200 55088 320000 55208 6 la_data_out[50]
port 319 nsew signal output
rlabel metal3 s 319200 56176 320000 56296 6 la_data_out[51]
port 320 nsew signal output
rlabel metal3 s 319200 57400 320000 57520 6 la_data_out[52]
port 321 nsew signal output
rlabel metal3 s 319200 58488 320000 58608 6 la_data_out[53]
port 322 nsew signal output
rlabel metal3 s 319200 59576 320000 59696 6 la_data_out[54]
port 323 nsew signal output
rlabel metal3 s 319200 60664 320000 60784 6 la_data_out[55]
port 324 nsew signal output
rlabel metal3 s 319200 61752 320000 61872 6 la_data_out[56]
port 325 nsew signal output
rlabel metal3 s 319200 62840 320000 62960 6 la_data_out[57]
port 326 nsew signal output
rlabel metal3 s 319200 63928 320000 64048 6 la_data_out[58]
port 327 nsew signal output
rlabel metal3 s 319200 65016 320000 65136 6 la_data_out[59]
port 328 nsew signal output
rlabel metal3 s 319200 5992 320000 6112 6 la_data_out[5]
port 329 nsew signal output
rlabel metal3 s 319200 66104 320000 66224 6 la_data_out[60]
port 330 nsew signal output
rlabel metal3 s 319200 67192 320000 67312 6 la_data_out[61]
port 331 nsew signal output
rlabel metal3 s 319200 68280 320000 68400 6 la_data_out[62]
port 332 nsew signal output
rlabel metal3 s 319200 69368 320000 69488 6 la_data_out[63]
port 333 nsew signal output
rlabel metal3 s 319200 70456 320000 70576 6 la_data_out[64]
port 334 nsew signal output
rlabel metal3 s 319200 71544 320000 71664 6 la_data_out[65]
port 335 nsew signal output
rlabel metal3 s 319200 72632 320000 72752 6 la_data_out[66]
port 336 nsew signal output
rlabel metal3 s 319200 73720 320000 73840 6 la_data_out[67]
port 337 nsew signal output
rlabel metal3 s 319200 74808 320000 74928 6 la_data_out[68]
port 338 nsew signal output
rlabel metal3 s 319200 75896 320000 76016 6 la_data_out[69]
port 339 nsew signal output
rlabel metal3 s 319200 7080 320000 7200 6 la_data_out[6]
port 340 nsew signal output
rlabel metal3 s 319200 76984 320000 77104 6 la_data_out[70]
port 341 nsew signal output
rlabel metal3 s 319200 78072 320000 78192 6 la_data_out[71]
port 342 nsew signal output
rlabel metal3 s 319200 79160 320000 79280 6 la_data_out[72]
port 343 nsew signal output
rlabel metal3 s 319200 80248 320000 80368 6 la_data_out[73]
port 344 nsew signal output
rlabel metal3 s 319200 81336 320000 81456 6 la_data_out[74]
port 345 nsew signal output
rlabel metal3 s 319200 82424 320000 82544 6 la_data_out[75]
port 346 nsew signal output
rlabel metal3 s 319200 83512 320000 83632 6 la_data_out[76]
port 347 nsew signal output
rlabel metal3 s 319200 84736 320000 84856 6 la_data_out[77]
port 348 nsew signal output
rlabel metal3 s 319200 85824 320000 85944 6 la_data_out[78]
port 349 nsew signal output
rlabel metal3 s 319200 86912 320000 87032 6 la_data_out[79]
port 350 nsew signal output
rlabel metal3 s 319200 8168 320000 8288 6 la_data_out[7]
port 351 nsew signal output
rlabel metal3 s 319200 88000 320000 88120 6 la_data_out[80]
port 352 nsew signal output
rlabel metal3 s 319200 89088 320000 89208 6 la_data_out[81]
port 353 nsew signal output
rlabel metal3 s 319200 90176 320000 90296 6 la_data_out[82]
port 354 nsew signal output
rlabel metal3 s 319200 91264 320000 91384 6 la_data_out[83]
port 355 nsew signal output
rlabel metal3 s 319200 92352 320000 92472 6 la_data_out[84]
port 356 nsew signal output
rlabel metal3 s 319200 93440 320000 93560 6 la_data_out[85]
port 357 nsew signal output
rlabel metal3 s 319200 94528 320000 94648 6 la_data_out[86]
port 358 nsew signal output
rlabel metal3 s 319200 95616 320000 95736 6 la_data_out[87]
port 359 nsew signal output
rlabel metal3 s 319200 96704 320000 96824 6 la_data_out[88]
port 360 nsew signal output
rlabel metal3 s 319200 97792 320000 97912 6 la_data_out[89]
port 361 nsew signal output
rlabel metal3 s 319200 9256 320000 9376 6 la_data_out[8]
port 362 nsew signal output
rlabel metal3 s 319200 98880 320000 99000 6 la_data_out[90]
port 363 nsew signal output
rlabel metal3 s 319200 99968 320000 100088 6 la_data_out[91]
port 364 nsew signal output
rlabel metal3 s 319200 101056 320000 101176 6 la_data_out[92]
port 365 nsew signal output
rlabel metal3 s 319200 102144 320000 102264 6 la_data_out[93]
port 366 nsew signal output
rlabel metal3 s 319200 103232 320000 103352 6 la_data_out[94]
port 367 nsew signal output
rlabel metal3 s 319200 104320 320000 104440 6 la_data_out[95]
port 368 nsew signal output
rlabel metal3 s 319200 105408 320000 105528 6 la_data_out[96]
port 369 nsew signal output
rlabel metal3 s 319200 106496 320000 106616 6 la_data_out[97]
port 370 nsew signal output
rlabel metal3 s 319200 107584 320000 107704 6 la_data_out[98]
port 371 nsew signal output
rlabel metal3 s 319200 108672 320000 108792 6 la_data_out[99]
port 372 nsew signal output
rlabel metal3 s 319200 10344 320000 10464 6 la_data_out[9]
port 373 nsew signal output
rlabel metal3 s 0 70184 800 70304 6 la_oenb[0]
port 374 nsew signal input
rlabel metal3 s 0 124856 800 124976 6 la_oenb[100]
port 375 nsew signal input
rlabel metal3 s 0 125400 800 125520 6 la_oenb[101]
port 376 nsew signal input
rlabel metal3 s 0 125944 800 126064 6 la_oenb[102]
port 377 nsew signal input
rlabel metal3 s 0 126488 800 126608 6 la_oenb[103]
port 378 nsew signal input
rlabel metal3 s 0 127032 800 127152 6 la_oenb[104]
port 379 nsew signal input
rlabel metal3 s 0 127576 800 127696 6 la_oenb[105]
port 380 nsew signal input
rlabel metal3 s 0 128120 800 128240 6 la_oenb[106]
port 381 nsew signal input
rlabel metal3 s 0 128664 800 128784 6 la_oenb[107]
port 382 nsew signal input
rlabel metal3 s 0 129208 800 129328 6 la_oenb[108]
port 383 nsew signal input
rlabel metal3 s 0 129752 800 129872 6 la_oenb[109]
port 384 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 la_oenb[10]
port 385 nsew signal input
rlabel metal3 s 0 130296 800 130416 6 la_oenb[110]
port 386 nsew signal input
rlabel metal3 s 0 130840 800 130960 6 la_oenb[111]
port 387 nsew signal input
rlabel metal3 s 0 131384 800 131504 6 la_oenb[112]
port 388 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 la_oenb[113]
port 389 nsew signal input
rlabel metal3 s 0 132472 800 132592 6 la_oenb[114]
port 390 nsew signal input
rlabel metal3 s 0 133016 800 133136 6 la_oenb[115]
port 391 nsew signal input
rlabel metal3 s 0 133560 800 133680 6 la_oenb[116]
port 392 nsew signal input
rlabel metal3 s 0 134104 800 134224 6 la_oenb[117]
port 393 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 la_oenb[118]
port 394 nsew signal input
rlabel metal3 s 0 135192 800 135312 6 la_oenb[119]
port 395 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 la_oenb[11]
port 396 nsew signal input
rlabel metal3 s 0 135736 800 135856 6 la_oenb[120]
port 397 nsew signal input
rlabel metal3 s 0 136280 800 136400 6 la_oenb[121]
port 398 nsew signal input
rlabel metal3 s 0 136824 800 136944 6 la_oenb[122]
port 399 nsew signal input
rlabel metal3 s 0 137368 800 137488 6 la_oenb[123]
port 400 nsew signal input
rlabel metal3 s 0 137912 800 138032 6 la_oenb[124]
port 401 nsew signal input
rlabel metal3 s 0 138456 800 138576 6 la_oenb[125]
port 402 nsew signal input
rlabel metal3 s 0 139000 800 139120 6 la_oenb[126]
port 403 nsew signal input
rlabel metal3 s 0 139544 800 139664 6 la_oenb[127]
port 404 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 la_oenb[12]
port 405 nsew signal input
rlabel metal3 s 0 77256 800 77376 6 la_oenb[13]
port 406 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 la_oenb[14]
port 407 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 la_oenb[15]
port 408 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 la_oenb[16]
port 409 nsew signal input
rlabel metal3 s 0 79432 800 79552 6 la_oenb[17]
port 410 nsew signal input
rlabel metal3 s 0 79976 800 80096 6 la_oenb[18]
port 411 nsew signal input
rlabel metal3 s 0 80520 800 80640 6 la_oenb[19]
port 412 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 la_oenb[1]
port 413 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 la_oenb[20]
port 414 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 la_oenb[21]
port 415 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 la_oenb[22]
port 416 nsew signal input
rlabel metal3 s 0 82696 800 82816 6 la_oenb[23]
port 417 nsew signal input
rlabel metal3 s 0 83240 800 83360 6 la_oenb[24]
port 418 nsew signal input
rlabel metal3 s 0 83784 800 83904 6 la_oenb[25]
port 419 nsew signal input
rlabel metal3 s 0 84464 800 84584 6 la_oenb[26]
port 420 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 la_oenb[27]
port 421 nsew signal input
rlabel metal3 s 0 85552 800 85672 6 la_oenb[28]
port 422 nsew signal input
rlabel metal3 s 0 86096 800 86216 6 la_oenb[29]
port 423 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 la_oenb[2]
port 424 nsew signal input
rlabel metal3 s 0 86640 800 86760 6 la_oenb[30]
port 425 nsew signal input
rlabel metal3 s 0 87184 800 87304 6 la_oenb[31]
port 426 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 la_oenb[32]
port 427 nsew signal input
rlabel metal3 s 0 88272 800 88392 6 la_oenb[33]
port 428 nsew signal input
rlabel metal3 s 0 88816 800 88936 6 la_oenb[34]
port 429 nsew signal input
rlabel metal3 s 0 89360 800 89480 6 la_oenb[35]
port 430 nsew signal input
rlabel metal3 s 0 89904 800 90024 6 la_oenb[36]
port 431 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 la_oenb[37]
port 432 nsew signal input
rlabel metal3 s 0 90992 800 91112 6 la_oenb[38]
port 433 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 la_oenb[39]
port 434 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 la_oenb[3]
port 435 nsew signal input
rlabel metal3 s 0 92080 800 92200 6 la_oenb[40]
port 436 nsew signal input
rlabel metal3 s 0 92624 800 92744 6 la_oenb[41]
port 437 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 la_oenb[42]
port 438 nsew signal input
rlabel metal3 s 0 93712 800 93832 6 la_oenb[43]
port 439 nsew signal input
rlabel metal3 s 0 94256 800 94376 6 la_oenb[44]
port 440 nsew signal input
rlabel metal3 s 0 94800 800 94920 6 la_oenb[45]
port 441 nsew signal input
rlabel metal3 s 0 95344 800 95464 6 la_oenb[46]
port 442 nsew signal input
rlabel metal3 s 0 95888 800 96008 6 la_oenb[47]
port 443 nsew signal input
rlabel metal3 s 0 96432 800 96552 6 la_oenb[48]
port 444 nsew signal input
rlabel metal3 s 0 96976 800 97096 6 la_oenb[49]
port 445 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 la_oenb[4]
port 446 nsew signal input
rlabel metal3 s 0 97520 800 97640 6 la_oenb[50]
port 447 nsew signal input
rlabel metal3 s 0 98064 800 98184 6 la_oenb[51]
port 448 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 la_oenb[52]
port 449 nsew signal input
rlabel metal3 s 0 99152 800 99272 6 la_oenb[53]
port 450 nsew signal input
rlabel metal3 s 0 99696 800 99816 6 la_oenb[54]
port 451 nsew signal input
rlabel metal3 s 0 100240 800 100360 6 la_oenb[55]
port 452 nsew signal input
rlabel metal3 s 0 100784 800 100904 6 la_oenb[56]
port 453 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 la_oenb[57]
port 454 nsew signal input
rlabel metal3 s 0 101872 800 101992 6 la_oenb[58]
port 455 nsew signal input
rlabel metal3 s 0 102416 800 102536 6 la_oenb[59]
port 456 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 la_oenb[5]
port 457 nsew signal input
rlabel metal3 s 0 102960 800 103080 6 la_oenb[60]
port 458 nsew signal input
rlabel metal3 s 0 103504 800 103624 6 la_oenb[61]
port 459 nsew signal input
rlabel metal3 s 0 104048 800 104168 6 la_oenb[62]
port 460 nsew signal input
rlabel metal3 s 0 104592 800 104712 6 la_oenb[63]
port 461 nsew signal input
rlabel metal3 s 0 105136 800 105256 6 la_oenb[64]
port 462 nsew signal input
rlabel metal3 s 0 105680 800 105800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal3 s 0 106224 800 106344 6 la_oenb[66]
port 464 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 la_oenb[67]
port 465 nsew signal input
rlabel metal3 s 0 107312 800 107432 6 la_oenb[68]
port 466 nsew signal input
rlabel metal3 s 0 107856 800 107976 6 la_oenb[69]
port 467 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 la_oenb[6]
port 468 nsew signal input
rlabel metal3 s 0 108400 800 108520 6 la_oenb[70]
port 469 nsew signal input
rlabel metal3 s 0 108944 800 109064 6 la_oenb[71]
port 470 nsew signal input
rlabel metal3 s 0 109488 800 109608 6 la_oenb[72]
port 471 nsew signal input
rlabel metal3 s 0 110032 800 110152 6 la_oenb[73]
port 472 nsew signal input
rlabel metal3 s 0 110576 800 110696 6 la_oenb[74]
port 473 nsew signal input
rlabel metal3 s 0 111120 800 111240 6 la_oenb[75]
port 474 nsew signal input
rlabel metal3 s 0 111664 800 111784 6 la_oenb[76]
port 475 nsew signal input
rlabel metal3 s 0 112344 800 112464 6 la_oenb[77]
port 476 nsew signal input
rlabel metal3 s 0 112888 800 113008 6 la_oenb[78]
port 477 nsew signal input
rlabel metal3 s 0 113432 800 113552 6 la_oenb[79]
port 478 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 la_oenb[7]
port 479 nsew signal input
rlabel metal3 s 0 113976 800 114096 6 la_oenb[80]
port 480 nsew signal input
rlabel metal3 s 0 114520 800 114640 6 la_oenb[81]
port 481 nsew signal input
rlabel metal3 s 0 115064 800 115184 6 la_oenb[82]
port 482 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 la_oenb[83]
port 483 nsew signal input
rlabel metal3 s 0 116152 800 116272 6 la_oenb[84]
port 484 nsew signal input
rlabel metal3 s 0 116696 800 116816 6 la_oenb[85]
port 485 nsew signal input
rlabel metal3 s 0 117240 800 117360 6 la_oenb[86]
port 486 nsew signal input
rlabel metal3 s 0 117784 800 117904 6 la_oenb[87]
port 487 nsew signal input
rlabel metal3 s 0 118328 800 118448 6 la_oenb[88]
port 488 nsew signal input
rlabel metal3 s 0 118872 800 118992 6 la_oenb[89]
port 489 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 la_oenb[8]
port 490 nsew signal input
rlabel metal3 s 0 119416 800 119536 6 la_oenb[90]
port 491 nsew signal input
rlabel metal3 s 0 119960 800 120080 6 la_oenb[91]
port 492 nsew signal input
rlabel metal3 s 0 120504 800 120624 6 la_oenb[92]
port 493 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 la_oenb[93]
port 494 nsew signal input
rlabel metal3 s 0 121592 800 121712 6 la_oenb[94]
port 495 nsew signal input
rlabel metal3 s 0 122136 800 122256 6 la_oenb[95]
port 496 nsew signal input
rlabel metal3 s 0 122680 800 122800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal3 s 0 123224 800 123344 6 la_oenb[97]
port 498 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 la_oenb[98]
port 499 nsew signal input
rlabel metal3 s 0 124312 800 124432 6 la_oenb[99]
port 500 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 24208 2128 24528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 44208 2128 44528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 64208 2128 64528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 84208 2128 84528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 104208 2128 104528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 124208 2128 124528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 144208 2128 144528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 164208 2128 164528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 184208 2128 184528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 204208 2128 204528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 224208 2128 224528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 244208 2128 244528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 264208 2128 264528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 284208 2128 284528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 304208 2128 304528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 14208 2128 14528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 34208 2128 34528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 54208 2128 54528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 74208 2128 74528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 94208 2128 94528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 114208 2128 114528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 134208 2128 134528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 154208 2128 154528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 174208 2128 174528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 194208 2128 194528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 214208 2128 214528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234208 2128 234528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 254208 2128 254528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 274208 2128 274528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 294208 2128 294528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 314208 2128 314528 137680 6 vssd1
port 503 nsew ground input
rlabel metal2 s 1398 0 1454 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 154026 0 154082 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 171598 0 171654 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 180430 0 180486 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 189262 0 189318 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 198002 0 198058 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 206834 0 206890 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 215666 0 215722 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 224498 0 224554 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 233238 0 233294 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 242070 0 242126 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 250902 0 250958 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 259642 0 259698 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 268474 0 268530 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 277306 0 277362 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 286138 0 286194 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 294878 0 294934 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 303710 0 303766 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 165710 0 165766 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 174542 0 174598 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 183374 0 183430 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 192206 0 192262 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 200946 0 201002 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 209778 0 209834 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 218610 0 218666 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 227350 0 227406 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 236182 0 236238 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 245014 0 245070 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 253846 0 253902 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 262586 0 262642 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 271418 0 271474 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 280250 0 280306 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 289082 0 289138 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 297822 0 297878 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 306654 0 306710 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 112902 0 112958 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 133418 0 133474 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 142250 0 142306 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 151082 0 151138 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 159914 0 159970 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 168654 0 168710 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 177486 0 177542 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 186318 0 186374 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 195058 0 195114 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 203890 0 203946 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 212722 0 212778 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 221554 0 221610 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 230294 0 230350 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 239126 0 239182 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 247958 0 248014 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 256790 0 256846 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 265530 0 265586 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 274362 0 274418 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 283194 0 283250 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 291934 0 291990 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 300766 0 300822 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 309598 0 309654 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 98182 0 98238 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 107014 0 107070 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 320000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 141201008
string GDS_FILE /home/serdar/Desktop/pwm/pwm_openmpw/openlane/pwm/runs/pwm/results/finishing/pwm_top.magic.gds
string GDS_START 1703952
<< end >>

